-- HW_QSYS.vhd

-- Generated using ACDS version 15.1 185

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity HW_QSYS is
	port (
		clk_125_clk                                  : in    std_logic                     := '0';             --             clk_125.clk
		clk_50_clk                                   : in    std_logic                     := '0';             --              clk_50.clk
		i2c_scl_export                               : out   std_logic;                                        --             i2c_scl.export
		i2c_sda_export                               : inout std_logic                     := '0';             --             i2c_sda.export
		key_export                                   : in    std_logic_vector(3 downto 0)  := (others => '0'); --                 key.export
		ledg_export                                  : out   std_logic_vector(7 downto 0);                     --                ledg.export
		ledr_export                                  : out   std_logic_vector(7 downto 0);                     --                ledr.export
		lpddr2_mem_ca                                : out   std_logic_vector(9 downto 0);                     --              lpddr2.mem_ca
		lpddr2_mem_ck                                : out   std_logic_vector(0 downto 0);                     --                    .mem_ck
		lpddr2_mem_ck_n                              : out   std_logic_vector(0 downto 0);                     --                    .mem_ck_n
		lpddr2_mem_cke                               : out   std_logic_vector(0 downto 0);                     --                    .mem_cke
		lpddr2_mem_cs_n                              : out   std_logic_vector(0 downto 0);                     --                    .mem_cs_n
		lpddr2_mem_dm                                : out   std_logic_vector(3 downto 0);                     --                    .mem_dm
		lpddr2_mem_dq                                : inout std_logic_vector(31 downto 0) := (others => '0'); --                    .mem_dq
		lpddr2_mem_dqs                               : inout std_logic_vector(3 downto 0)  := (others => '0'); --                    .mem_dqs
		lpddr2_mem_dqs_n                             : inout std_logic_vector(3 downto 0)  := (others => '0'); --                    .mem_dqs_n
		lpddr2_global_reset_reset_n                  : in    std_logic                     := '0';             -- lpddr2_global_reset.reset_n
		lpddr2_oct_rzqin                             : in    std_logic                     := '0';             --          lpddr2_oct.rzqin
		lpddr2_pll_ref_clk_clk                       : in    std_logic                     := '0';             --  lpddr2_pll_ref_clk.clk
		lpddr2_pll_sharing_pll_mem_clk               : out   std_logic;                                        --  lpddr2_pll_sharing.pll_mem_clk
		lpddr2_pll_sharing_pll_write_clk             : out   std_logic;                                        --                    .pll_write_clk
		lpddr2_pll_sharing_pll_locked                : out   std_logic;                                        --                    .pll_locked
		lpddr2_pll_sharing_pll_write_clk_pre_phy_clk : out   std_logic;                                        --                    .pll_write_clk_pre_phy_clk
		lpddr2_pll_sharing_pll_addr_cmd_clk          : out   std_logic;                                        --                    .pll_addr_cmd_clk
		lpddr2_pll_sharing_pll_avl_clk               : out   std_logic;                                        --                    .pll_avl_clk
		lpddr2_pll_sharing_pll_config_clk            : out   std_logic;                                        --                    .pll_config_clk
		lpddr2_pll_sharing_pll_mem_phy_clk           : out   std_logic;                                        --                    .pll_mem_phy_clk
		lpddr2_pll_sharing_afi_phy_clk               : out   std_logic;                                        --                    .afi_phy_clk
		lpddr2_pll_sharing_pll_avl_phy_clk           : out   std_logic;                                        --                    .pll_avl_phy_clk
		lpddr2_status_local_init_done                : out   std_logic;                                        --       lpddr2_status.local_init_done
		lpddr2_status_local_cal_success              : out   std_logic;                                        --                    .local_cal_success
		lpddr2_status_local_cal_fail                 : out   std_logic;                                        --                    .local_cal_fail
		reset_reset_n                                : in    std_logic                     := '0';             --               reset.reset_n
		sd_sd_clk                                    : out   std_logic;                                        --                  sd.sd_clk
		sd_sd_cmd                                    : inout std_logic                     := '0';             --                    .sd_cmd
		sd_sd_dat                                    : inout std_logic_vector(3 downto 0)  := (others => '0'); --                    .sd_dat
		sram_bridge_out_sram_tcm_data_out            : inout std_logic_vector(15 downto 0) := (others => '0'); --     sram_bridge_out.sram_tcm_data_out
		sram_bridge_out_sram_tcm_address_out         : out   std_logic_vector(18 downto 0);                    --                    .sram_tcm_address_out
		sram_bridge_out_sram_tcm_outputenable_n_out  : out   std_logic_vector(0 downto 0);                     --                    .sram_tcm_outputenable_n_out
		sram_bridge_out_sram_tcm_chipselect_n_out    : out   std_logic_vector(0 downto 0);                     --                    .sram_tcm_chipselect_n_out
		sram_bridge_out_sram_tcm_byteenable_n_out    : out   std_logic_vector(1 downto 0);                     --                    .sram_tcm_byteenable_n_out
		sram_bridge_out_sram_tcm_write_n_out         : out   std_logic_vector(0 downto 0);                     --                    .sram_tcm_write_n_out
		video_RGB_OUT                                : out   std_logic_vector(23 downto 0);                    --               video.RGB_OUT
		video_HD                                     : out   std_logic;                                        --                    .HD
		video_VD                                     : out   std_logic;                                        --                    .VD
		video_DEN                                    : out   std_logic;                                        --                    .DEN
		video_clk_clk                                : out   std_logic                                         --           video_clk.clk
	);
end entity HW_QSYS;

architecture rtl of HW_QSYS is
	component Pixel_Conv is
		generic (
			SOURCE_SYMBOLS_PER_BEAT : integer := 3
		);
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			reset_n   : in  std_logic                     := 'X';             -- reset_n
			ready_out : out std_logic;                                        -- ready
			valid_in  : in  std_logic                     := 'X';             -- valid
			data_in   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			eop_in    : in  std_logic                     := 'X';             -- endofpacket
			sop_in    : in  std_logic                     := 'X';             -- startofpacket
			empty_in  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			ready_in  : in  std_logic                     := 'X';             -- ready
			valid_out : out std_logic;                                        -- valid
			data_out  : out std_logic_vector(23 downto 0);                    -- data
			eop_out   : out std_logic;                                        -- endofpacket
			sop_out   : out std_logic;                                        -- startofpacket
			empty_out : out std_logic                                         -- empty
		);
	end component Pixel_Conv;

	component HW_QSYS_cpu_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(29 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_burstcount                        : out std_logic_vector(3 downto 0);                     -- burstcount
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(29 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component HW_QSYS_cpu_0;

	component HW_QSYS_cpu_1 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(29 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_burstcount                        : out std_logic_vector(3 downto 0);                     -- burstcount
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(29 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component HW_QSYS_cpu_1;

	component HW_QSYS_cpu_2 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(29 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_burstcount                        : out std_logic_vector(3 downto 0);                     -- burstcount
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(29 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component HW_QSYS_cpu_2;

	component HW_QSYS_i2c_scl is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component HW_QSYS_i2c_scl;

	component HW_QSYS_i2c_sda is
		port (
			clk        : in    std_logic                     := 'X';             -- clk
			reset_n    : in    std_logic                     := 'X';             -- reset_n
			address    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in    std_logic                     := 'X';             -- write_n
			writedata  : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in    std_logic                     := 'X';             -- chipselect
			readdata   : out   std_logic_vector(31 downto 0);                    -- readdata
			bidir_port : inout std_logic                     := 'X'              -- export
		);
	end component HW_QSYS_i2c_sda;

	component HW_QSYS_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component HW_QSYS_jtag_uart_0;

	component HW_QSYS_key is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component HW_QSYS_key;

	component HW_QSYS_ledg is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component HW_QSYS_ledg;

	component HW_QSYS_lpddr2 is
		port (
			pll_ref_clk                : in    std_logic                     := 'X';             -- clk
			global_reset_n             : in    std_logic                     := 'X';             -- reset_n
			soft_reset_n               : in    std_logic                     := 'X';             -- reset_n
			afi_clk                    : out   std_logic;                                        -- clk
			afi_half_clk               : out   std_logic;                                        -- clk
			afi_reset_n                : out   std_logic;                                        -- reset_n
			afi_reset_export_n         : out   std_logic;                                        -- reset_n
			mem_ca                     : out   std_logic_vector(9 downto 0);                     -- mem_ca
			mem_ck                     : out   std_logic_vector(0 downto 0);                     -- mem_ck
			mem_ck_n                   : out   std_logic_vector(0 downto 0);                     -- mem_ck_n
			mem_cke                    : out   std_logic_vector(0 downto 0);                     -- mem_cke
			mem_cs_n                   : out   std_logic_vector(0 downto 0);                     -- mem_cs_n
			mem_dm                     : out   std_logic_vector(3 downto 0);                     -- mem_dm
			mem_dq                     : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs                    : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n                  : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
			avl_ready_0                : out   std_logic;                                        -- waitrequest_n
			avl_burstbegin_0           : in    std_logic                     := 'X';             -- beginbursttransfer
			avl_addr_0                 : in    std_logic_vector(26 downto 0) := (others => 'X'); -- address
			avl_rdata_valid_0          : out   std_logic;                                        -- readdatavalid
			avl_rdata_0                : out   std_logic_vector(31 downto 0);                    -- readdata
			avl_wdata_0                : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avl_be_0                   : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avl_read_req_0             : in    std_logic                     := 'X';             -- read
			avl_write_req_0            : in    std_logic                     := 'X';             -- write
			avl_size_0                 : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- burstcount
			avl_ready_1                : out   std_logic;                                        -- waitrequest_n
			avl_burstbegin_1           : in    std_logic                     := 'X';             -- beginbursttransfer
			avl_addr_1                 : in    std_logic_vector(26 downto 0) := (others => 'X'); -- address
			avl_rdata_valid_1          : out   std_logic;                                        -- readdatavalid
			avl_rdata_1                : out   std_logic_vector(31 downto 0);                    -- readdata
			avl_wdata_1                : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avl_be_1                   : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avl_read_req_1             : in    std_logic                     := 'X';             -- read
			avl_write_req_1            : in    std_logic                     := 'X';             -- write
			avl_size_1                 : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- burstcount
			avl_ready_2                : out   std_logic;                                        -- waitrequest_n
			avl_burstbegin_2           : in    std_logic                     := 'X';             -- beginbursttransfer
			avl_addr_2                 : in    std_logic_vector(26 downto 0) := (others => 'X'); -- address
			avl_rdata_valid_2          : out   std_logic;                                        -- readdatavalid
			avl_rdata_2                : out   std_logic_vector(31 downto 0);                    -- readdata
			avl_wdata_2                : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avl_be_2                   : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avl_read_req_2             : in    std_logic                     := 'X';             -- read
			avl_write_req_2            : in    std_logic                     := 'X';             -- write
			avl_size_2                 : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- burstcount
			mp_cmd_clk_0_clk           : in    std_logic                     := 'X';             -- clk
			mp_cmd_reset_n_0_reset_n   : in    std_logic                     := 'X';             -- reset_n
			mp_cmd_clk_1_clk           : in    std_logic                     := 'X';             -- clk
			mp_cmd_reset_n_1_reset_n   : in    std_logic                     := 'X';             -- reset_n
			mp_cmd_clk_2_clk           : in    std_logic                     := 'X';             -- clk
			mp_cmd_reset_n_2_reset_n   : in    std_logic                     := 'X';             -- reset_n
			mp_rfifo_clk_0_clk         : in    std_logic                     := 'X';             -- clk
			mp_rfifo_reset_n_0_reset_n : in    std_logic                     := 'X';             -- reset_n
			mp_wfifo_clk_0_clk         : in    std_logic                     := 'X';             -- clk
			mp_wfifo_reset_n_0_reset_n : in    std_logic                     := 'X';             -- reset_n
			mp_rfifo_clk_1_clk         : in    std_logic                     := 'X';             -- clk
			mp_rfifo_reset_n_1_reset_n : in    std_logic                     := 'X';             -- reset_n
			mp_wfifo_clk_1_clk         : in    std_logic                     := 'X';             -- clk
			mp_wfifo_reset_n_1_reset_n : in    std_logic                     := 'X';             -- reset_n
			local_init_done            : out   std_logic;                                        -- local_init_done
			local_cal_success          : out   std_logic;                                        -- local_cal_success
			local_cal_fail             : out   std_logic;                                        -- local_cal_fail
			oct_rzqin                  : in    std_logic                     := 'X';             -- rzqin
			pll_mem_clk                : out   std_logic;                                        -- pll_mem_clk
			pll_write_clk              : out   std_logic;                                        -- pll_write_clk
			pll_locked                 : out   std_logic;                                        -- pll_locked
			pll_write_clk_pre_phy_clk  : out   std_logic;                                        -- pll_write_clk_pre_phy_clk
			pll_addr_cmd_clk           : out   std_logic;                                        -- pll_addr_cmd_clk
			pll_avl_clk                : out   std_logic;                                        -- pll_avl_clk
			pll_config_clk             : out   std_logic;                                        -- pll_config_clk
			pll_mem_phy_clk            : out   std_logic;                                        -- pll_mem_phy_clk
			afi_phy_clk                : out   std_logic;                                        -- afi_phy_clk
			pll_avl_phy_clk            : out   std_logic                                         -- pll_avl_phy_clk
		);
	end component HW_QSYS_lpddr2;

	component altera_avalon_mailbox is
		generic (
			DWIDTH : integer := 32;
			AWIDTH : integer := 2
		);
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			rst_n                : in  std_logic                     := 'X';             -- reset_n
			avmm_snd_address     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			avmm_snd_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avmm_snd_write       : in  std_logic                     := 'X';             -- write
			avmm_snd_read        : in  std_logic                     := 'X';             -- read
			avmm_snd_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			avmm_snd_waitrequest : out std_logic;                                        -- waitrequest
			irq_msg              : out std_logic;                                        -- irq
			avmm_rcv_address     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			avmm_rcv_read        : in  std_logic                     := 'X';             -- read
			avmm_rcv_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avmm_rcv_write       : in  std_logic                     := 'X';             -- write
			avmm_rcv_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			irq_space            : out std_logic                                         -- irq
		);
	end component altera_avalon_mailbox;

	component HW_QSYS_read_dma_0 is
		port (
			mm_read_address              : out std_logic_vector(28 downto 0);                     -- address
			mm_read_read                 : out std_logic;                                         -- read
			mm_read_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			mm_read_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			mm_read_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			mm_read_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			mm_read_burstcount           : out std_logic_vector(7 downto 0);                      -- burstcount
			clock_clk                    : in  std_logic                      := 'X';             -- clk
			reset_n_reset_n              : in  std_logic                      := 'X';             -- reset_n
			csr_writedata                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			csr_write                    : in  std_logic                      := 'X';             -- write
			csr_byteenable               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			csr_readdata                 : out std_logic_vector(31 downto 0);                     -- readdata
			csr_read                     : in  std_logic                      := 'X';             -- read
			csr_address                  : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- address
			descriptor_slave_write       : in  std_logic                      := 'X';             -- write
			descriptor_slave_waitrequest : out std_logic;                                         -- waitrequest
			descriptor_slave_writedata   : in  std_logic_vector(127 downto 0) := (others => 'X'); -- writedata
			descriptor_slave_byteenable  : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- byteenable
			csr_irq_irq                  : out std_logic;                                         -- irq
			st_source_data               : out std_logic_vector(31 downto 0);                     -- data
			st_source_valid              : out std_logic;                                         -- valid
			st_source_ready              : in  std_logic                      := 'X'              -- ready
		);
	end component HW_QSYS_read_dma_0;

	component sd_cont is
		port (
			clk             : in    std_logic                     := 'X';             -- clk
			reset           : in    std_logic                     := 'X';             -- reset
			s_address       : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			s_read          : in    std_logic                     := 'X';             -- read
			s_readdata      : out   std_logic_vector(31 downto 0);                    -- readdata
			s_write         : in    std_logic                     := 'X';             -- write
			s_writedata     : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s_chipselect    : in    std_logic                     := 'X';             -- chipselect
			s_waitrequest_n : out   std_logic;                                        -- waitrequest_n
			m_address       : out   std_logic_vector(31 downto 0);                    -- address
			m_read          : out   std_logic;                                        -- read
			m_readdata      : in    std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m_write         : out   std_logic;                                        -- write
			m_writedata     : out   std_logic_vector(31 downto 0);                    -- writedata
			m_waitrequest_n : in    std_logic                     := 'X';             -- waitrequest_n
			sd_clk          : out   std_logic;                                        -- sd_clk
			sd_cmd          : inout std_logic                     := 'X';             -- sd_cmd
			sd_dat          : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- sd_dat
			sd_pll_clk      : in    std_logic                     := 'X'              -- clk
		);
	end component sd_cont;

	component HW_QSYS_sram is
		generic (
			TCM_ADDRESS_W                  : integer := 30;
			TCM_DATA_W                     : integer := 32;
			TCM_BYTEENABLE_W               : integer := 4;
			TCM_READ_WAIT                  : integer := 1;
			TCM_WRITE_WAIT                 : integer := 0;
			TCM_SETUP_WAIT                 : integer := 0;
			TCM_DATA_HOLD                  : integer := 0;
			TCM_TURNAROUND_TIME            : integer := 2;
			TCM_TIMING_UNITS               : integer := 1;
			TCM_READLATENCY                : integer := 2;
			TCM_SYMBOLS_PER_WORD           : integer := 4;
			USE_READDATA                   : integer := 1;
			USE_WRITEDATA                  : integer := 1;
			USE_READ                       : integer := 1;
			USE_WRITE                      : integer := 1;
			USE_BYTEENABLE                 : integer := 1;
			USE_CHIPSELECT                 : integer := 0;
			USE_LOCK                       : integer := 0;
			USE_ADDRESS                    : integer := 1;
			USE_WAITREQUEST                : integer := 0;
			USE_WRITEBYTEENABLE            : integer := 0;
			USE_OUTPUTENABLE               : integer := 0;
			USE_RESETREQUEST               : integer := 0;
			USE_IRQ                        : integer := 0;
			USE_RESET_OUTPUT               : integer := 0;
			ACTIVE_LOW_READ                : integer := 0;
			ACTIVE_LOW_LOCK                : integer := 0;
			ACTIVE_LOW_WRITE               : integer := 0;
			ACTIVE_LOW_CHIPSELECT          : integer := 0;
			ACTIVE_LOW_BYTEENABLE          : integer := 0;
			ACTIVE_LOW_OUTPUTENABLE        : integer := 0;
			ACTIVE_LOW_WRITEBYTEENABLE     : integer := 0;
			ACTIVE_LOW_WAITREQUEST         : integer := 0;
			ACTIVE_LOW_BEGINTRANSFER       : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0
		);
		port (
			clk_clk                : in  std_logic                     := 'X';             -- clk
			reset_reset            : in  std_logic                     := 'X';             -- reset
			uas_address            : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			uas_burstcount         : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- burstcount
			uas_read               : in  std_logic                     := 'X';             -- read
			uas_write              : in  std_logic                     := 'X';             -- write
			uas_waitrequest        : out std_logic;                                        -- waitrequest
			uas_readdatavalid      : out std_logic;                                        -- readdatavalid
			uas_byteenable         : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			uas_readdata           : out std_logic_vector(15 downto 0);                    -- readdata
			uas_writedata          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			uas_lock               : in  std_logic                     := 'X';             -- lock
			uas_debugaccess        : in  std_logic                     := 'X';             -- debugaccess
			tcm_write_n_out        : out std_logic;                                        -- write_n_out
			tcm_chipselect_n_out   : out std_logic;                                        -- chipselect_n_out
			tcm_outputenable_n_out : out std_logic;                                        -- outputenable_n_out
			tcm_request            : out std_logic;                                        -- request
			tcm_grant              : in  std_logic                     := 'X';             -- grant
			tcm_address_out        : out std_logic_vector(18 downto 0);                    -- address_out
			tcm_byteenable_n_out   : out std_logic_vector(1 downto 0);                     -- byteenable_n_out
			tcm_data_out           : out std_logic_vector(15 downto 0);                    -- data_out
			tcm_data_outen         : out std_logic;                                        -- data_outen
			tcm_data_in            : in  std_logic_vector(15 downto 0) := (others => 'X')  -- data_in
		);
	end component HW_QSYS_sram;

	component HW_QSYS_sram_bridge is
		port (
			clk                             : in    std_logic                     := 'X';             -- clk
			reset                           : in    std_logic                     := 'X';             -- reset
			request                         : in    std_logic                     := 'X';             -- request
			grant                           : out   std_logic;                                        -- grant
			tcs_sram_tcm_data_out           : in    std_logic_vector(15 downto 0) := (others => 'X'); -- sram_tcm_data_out_out
			tcs_sram_tcm_data_outen         : in    std_logic                     := 'X';             -- sram_tcm_data_out_outen
			tcs_sram_tcm_data_in            : out   std_logic_vector(15 downto 0);                    -- sram_tcm_data_out_in
			tcs_sram_tcm_address_out        : in    std_logic_vector(18 downto 0) := (others => 'X'); -- sram_tcm_address_out_out
			tcs_sram_tcm_outputenable_n_out : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- sram_tcm_outputenable_n_out_out
			tcs_sram_tcm_chipselect_n_out   : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- sram_tcm_chipselect_n_out_out
			tcs_sram_tcm_byteenable_n_out   : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- sram_tcm_byteenable_n_out_out
			tcs_sram_tcm_write_n_out        : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- sram_tcm_write_n_out_out
			sram_tcm_data_out               : inout std_logic_vector(15 downto 0) := (others => 'X'); -- sram_tcm_data_out
			sram_tcm_address_out            : out   std_logic_vector(18 downto 0);                    -- sram_tcm_address_out
			sram_tcm_outputenable_n_out     : out   std_logic_vector(0 downto 0);                     -- sram_tcm_outputenable_n_out
			sram_tcm_chipselect_n_out       : out   std_logic_vector(0 downto 0);                     -- sram_tcm_chipselect_n_out
			sram_tcm_byteenable_n_out       : out   std_logic_vector(1 downto 0);                     -- sram_tcm_byteenable_n_out
			sram_tcm_write_n_out            : out   std_logic_vector(0 downto 0)                      -- sram_tcm_write_n_out
		);
	end component HW_QSYS_sram_bridge;

	component HW_QSYS_sram_sharer is
		port (
			clk_clk                     : in  std_logic                     := 'X';             -- clk
			reset_reset                 : in  std_logic                     := 'X';             -- reset
			request                     : out std_logic;                                        -- request
			grant                       : in  std_logic                     := 'X';             -- grant
			sram_tcm_address_out        : out std_logic_vector(18 downto 0);                    -- sram_tcm_address_out_out
			sram_tcm_byteenable_n_out   : out std_logic_vector(1 downto 0);                     -- sram_tcm_byteenable_n_out_out
			sram_tcm_outputenable_n_out : out std_logic_vector(0 downto 0);                     -- sram_tcm_outputenable_n_out_out
			sram_tcm_write_n_out        : out std_logic_vector(0 downto 0);                     -- sram_tcm_write_n_out_out
			sram_tcm_data_out           : out std_logic_vector(15 downto 0);                    -- sram_tcm_data_out_out
			sram_tcm_data_in            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- sram_tcm_data_out_in
			sram_tcm_data_outen         : out std_logic;                                        -- sram_tcm_data_out_outen
			sram_tcm_chipselect_n_out   : out std_logic_vector(0 downto 0);                     -- sram_tcm_chipselect_n_out_out
			tcs0_request                : in  std_logic                     := 'X';             -- request
			tcs0_grant                  : out std_logic;                                        -- grant
			tcs0_address_out            : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address_out
			tcs0_byteenable_n_out       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n_out
			tcs0_outputenable_n_out     : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- outputenable_n_out
			tcs0_write_n_out            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- write_n_out
			tcs0_data_out               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data_out
			tcs0_data_in                : out std_logic_vector(15 downto 0);                    -- data_in
			tcs0_data_outen             : in  std_logic                     := 'X';             -- data_outen
			tcs0_chipselect_n_out       : in  std_logic_vector(0 downto 0)  := (others => 'X')  -- chipselect_n_out
		);
	end component HW_QSYS_sram_sharer;

	component HW_QSYS_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component HW_QSYS_sysid;

	component HW_QSYS_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component HW_QSYS_timer_0;

	component HW_QSYS_timer_1 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component HW_QSYS_timer_1;

	component twod_idct_st_hw is
		port (
			CLOCK     : in  std_logic                     := 'X';             -- clk
			DATAOUT   : out std_logic_vector(31 downto 0);                    -- data
			dst_ready : in  std_logic                     := 'X';             -- ready
			dst_valid : out std_logic;                                        -- valid
			reset     : in  std_logic                     := 'X';             -- reset
			DATAIN    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			src_ready : out std_logic;                                        -- ready
			src_valid : in  std_logic                     := 'X'              -- valid
		);
	end component twod_idct_st_hw;

	component altera_avalon_video_sync_generator is
		generic (
			DATA_STREAM_BIT_WIDTH : integer := 8;
			BEATS_PER_PIXEL       : integer := 3;
			NUM_COLUMNS           : integer := 800;
			NUM_ROWS              : integer := 480;
			H_BLANK_PIXELS        : integer := 216;
			H_FRONT_PORCH_PIXELS  : integer := 40;
			H_SYNC_PULSE_PIXELS   : integer := 1;
			H_SYNC_PULSE_POLARITY : integer := 0;
			V_BLANK_LINES         : integer := 35;
			V_FRONT_PORCH_LINES   : integer := 10;
			V_SYNC_PULSE_LINES    : integer := 1;
			V_SYNC_PULSE_POLARITY : integer := 0;
			TOTAL_HSCAN_PIXELS    : integer := 1056;
			TOTAL_VSCAN_LINES     : integer := 525
		);
		port (
			clk     : in  std_logic                     := 'X';             -- clk
			reset_n : in  std_logic                     := 'X';             -- reset_n
			ready   : out std_logic;                                        -- ready
			valid   : in  std_logic                     := 'X';             -- valid
			data    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			eop     : in  std_logic                     := 'X';             -- endofpacket
			sop     : in  std_logic                     := 'X';             -- startofpacket
			empty   : in  std_logic                     := 'X';             -- empty
			RGB_OUT : out std_logic_vector(23 downto 0);                    -- export
			HD      : out std_logic;                                        -- export
			VD      : out std_logic;                                        -- export
			DEN     : out std_logic                                         -- export
		);
	end component altera_avalon_video_sync_generator;

	component HW_QSYS_video_dma is
		port (
			mm_read_address              : out std_logic_vector(28 downto 0);                     -- address
			mm_read_read                 : out std_logic;                                         -- read
			mm_read_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			mm_read_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			mm_read_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			mm_read_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			mm_read_burstcount           : out std_logic_vector(7 downto 0);                      -- burstcount
			clock_clk                    : in  std_logic                      := 'X';             -- clk
			reset_n_reset_n              : in  std_logic                      := 'X';             -- reset_n
			csr_writedata                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			csr_write                    : in  std_logic                      := 'X';             -- write
			csr_byteenable               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			csr_readdata                 : out std_logic_vector(31 downto 0);                     -- readdata
			csr_read                     : in  std_logic                      := 'X';             -- read
			csr_address                  : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- address
			descriptor_slave_write       : in  std_logic                      := 'X';             -- write
			descriptor_slave_waitrequest : out std_logic;                                         -- waitrequest
			descriptor_slave_writedata   : in  std_logic_vector(127 downto 0) := (others => 'X'); -- writedata
			descriptor_slave_byteenable  : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- byteenable
			csr_irq_irq                  : out std_logic;                                         -- irq
			st_source_data               : out std_logic_vector(31 downto 0);                     -- data
			st_source_valid              : out std_logic;                                         -- valid
			st_source_ready              : in  std_logic                      := 'X';             -- ready
			st_source_startofpacket      : out std_logic;                                         -- startofpacket
			st_source_endofpacket        : out std_logic;                                         -- endofpacket
			st_source_empty              : out std_logic_vector(1 downto 0)                       -- empty
		);
	end component HW_QSYS_video_dma;

	component HW_QSYS_video_fifo is
		port (
			wrclock                       : in  std_logic                     := 'X';             -- clk
			wrreset_n                     : in  std_logic                     := 'X';             -- reset_n
			rdclock                       : in  std_logic                     := 'X';             -- clk
			rdreset_n                     : in  std_logic                     := 'X';             -- reset_n
			avalonst_sink_valid           : in  std_logic                     := 'X';             -- valid
			avalonst_sink_data            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			avalonst_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			avalonst_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			avalonst_sink_empty           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			avalonst_sink_ready           : out std_logic;                                        -- ready
			avalonst_source_valid         : out std_logic;                                        -- valid
			avalonst_source_data          : out std_logic_vector(31 downto 0);                    -- data
			avalonst_source_startofpacket : out std_logic;                                        -- startofpacket
			avalonst_source_endofpacket   : out std_logic;                                        -- endofpacket
			avalonst_source_empty         : out std_logic_vector(1 downto 0);                     -- empty
			avalonst_source_ready         : in  std_logic                     := 'X'              -- ready
		);
	end component HW_QSYS_video_fifo;

	component HW_QSYS_video_pll is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component HW_QSYS_video_pll;

	component HW_QSYS_write_dma_0 is
		port (
			mm_write_address             : out std_logic_vector(28 downto 0);                     -- address
			mm_write_write               : out std_logic;                                         -- write
			mm_write_byteenable          : out std_logic_vector(3 downto 0);                      -- byteenable
			mm_write_writedata           : out std_logic_vector(31 downto 0);                     -- writedata
			mm_write_waitrequest         : in  std_logic                      := 'X';             -- waitrequest
			mm_write_burstcount          : out std_logic_vector(7 downto 0);                      -- burstcount
			clock_clk                    : in  std_logic                      := 'X';             -- clk
			reset_n_reset_n              : in  std_logic                      := 'X';             -- reset_n
			csr_writedata                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			csr_write                    : in  std_logic                      := 'X';             -- write
			csr_byteenable               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			csr_readdata                 : out std_logic_vector(31 downto 0);                     -- readdata
			csr_read                     : in  std_logic                      := 'X';             -- read
			csr_address                  : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- address
			descriptor_slave_write       : in  std_logic                      := 'X';             -- write
			descriptor_slave_waitrequest : out std_logic;                                         -- waitrequest
			descriptor_slave_writedata   : in  std_logic_vector(127 downto 0) := (others => 'X'); -- writedata
			descriptor_slave_byteenable  : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- byteenable
			csr_irq_irq                  : out std_logic;                                         -- irq
			st_sink_data                 : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- data
			st_sink_valid                : in  std_logic                      := 'X';             -- valid
			st_sink_ready                : out std_logic                                          -- ready
		);
	end component HW_QSYS_write_dma_0;

	component HW_QSYS_mm_interconnect_0 is
		port (
			clk_125_clk_clk                                     : in  std_logic                      := 'X';             -- clk
			clk_50_out_clk_clk                                  : in  std_logic                      := 'X';             -- clk
			cpu_0_reset_reset_bridge_in_reset_reset             : in  std_logic                      := 'X';             -- reset
			cpu_1_reset_reset_bridge_in_reset_reset             : in  std_logic                      := 'X';             -- reset
			cpu_2_reset_reset_bridge_in_reset_reset             : in  std_logic                      := 'X';             -- reset
			lpddr2_mp_cmd_reset_n_0_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			mailbox_simple_1_rst_n_reset_bridge_in_reset_reset  : in  std_logic                      := 'X';             -- reset
			sd_cont_0_reset_reset_bridge_in_reset_reset         : in  std_logic                      := 'X';             -- reset
			cpu_0_data_master_address                           : in  std_logic_vector(29 downto 0)  := (others => 'X'); -- address
			cpu_0_data_master_waitrequest                       : out std_logic;                                         -- waitrequest
			cpu_0_data_master_burstcount                        : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- burstcount
			cpu_0_data_master_byteenable                        : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			cpu_0_data_master_read                              : in  std_logic                      := 'X';             -- read
			cpu_0_data_master_readdata                          : out std_logic_vector(31 downto 0);                     -- readdata
			cpu_0_data_master_readdatavalid                     : out std_logic;                                         -- readdatavalid
			cpu_0_data_master_write                             : in  std_logic                      := 'X';             -- write
			cpu_0_data_master_writedata                         : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			cpu_0_data_master_debugaccess                       : in  std_logic                      := 'X';             -- debugaccess
			cpu_0_instruction_master_address                    : in  std_logic_vector(29 downto 0)  := (others => 'X'); -- address
			cpu_0_instruction_master_waitrequest                : out std_logic;                                         -- waitrequest
			cpu_0_instruction_master_read                       : in  std_logic                      := 'X';             -- read
			cpu_0_instruction_master_readdata                   : out std_logic_vector(31 downto 0);                     -- readdata
			cpu_0_instruction_master_readdatavalid              : out std_logic;                                         -- readdatavalid
			cpu_1_data_master_address                           : in  std_logic_vector(29 downto 0)  := (others => 'X'); -- address
			cpu_1_data_master_waitrequest                       : out std_logic;                                         -- waitrequest
			cpu_1_data_master_burstcount                        : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- burstcount
			cpu_1_data_master_byteenable                        : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			cpu_1_data_master_read                              : in  std_logic                      := 'X';             -- read
			cpu_1_data_master_readdata                          : out std_logic_vector(31 downto 0);                     -- readdata
			cpu_1_data_master_readdatavalid                     : out std_logic;                                         -- readdatavalid
			cpu_1_data_master_write                             : in  std_logic                      := 'X';             -- write
			cpu_1_data_master_writedata                         : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			cpu_1_data_master_debugaccess                       : in  std_logic                      := 'X';             -- debugaccess
			cpu_1_instruction_master_address                    : in  std_logic_vector(29 downto 0)  := (others => 'X'); -- address
			cpu_1_instruction_master_waitrequest                : out std_logic;                                         -- waitrequest
			cpu_1_instruction_master_read                       : in  std_logic                      := 'X';             -- read
			cpu_1_instruction_master_readdata                   : out std_logic_vector(31 downto 0);                     -- readdata
			cpu_1_instruction_master_readdatavalid              : out std_logic;                                         -- readdatavalid
			cpu_2_data_master_address                           : in  std_logic_vector(29 downto 0)  := (others => 'X'); -- address
			cpu_2_data_master_waitrequest                       : out std_logic;                                         -- waitrequest
			cpu_2_data_master_burstcount                        : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- burstcount
			cpu_2_data_master_byteenable                        : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			cpu_2_data_master_read                              : in  std_logic                      := 'X';             -- read
			cpu_2_data_master_readdata                          : out std_logic_vector(31 downto 0);                     -- readdata
			cpu_2_data_master_readdatavalid                     : out std_logic;                                         -- readdatavalid
			cpu_2_data_master_write                             : in  std_logic                      := 'X';             -- write
			cpu_2_data_master_writedata                         : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			cpu_2_data_master_debugaccess                       : in  std_logic                      := 'X';             -- debugaccess
			cpu_2_instruction_master_address                    : in  std_logic_vector(29 downto 0)  := (others => 'X'); -- address
			cpu_2_instruction_master_waitrequest                : out std_logic;                                         -- waitrequest
			cpu_2_instruction_master_read                       : in  std_logic                      := 'X';             -- read
			cpu_2_instruction_master_readdata                   : out std_logic_vector(31 downto 0);                     -- readdata
			cpu_2_instruction_master_readdatavalid              : out std_logic;                                         -- readdatavalid
			sd_cont_0_master_address                            : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			sd_cont_0_master_waitrequest                        : out std_logic;                                         -- waitrequest
			sd_cont_0_master_read                               : in  std_logic                      := 'X';             -- read
			sd_cont_0_master_readdata                           : out std_logic_vector(31 downto 0);                     -- readdata
			sd_cont_0_master_write                              : in  std_logic                      := 'X';             -- write
			sd_cont_0_master_writedata                          : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			cpu_0_debug_mem_slave_address                       : out std_logic_vector(8 downto 0);                      -- address
			cpu_0_debug_mem_slave_write                         : out std_logic;                                         -- write
			cpu_0_debug_mem_slave_read                          : out std_logic;                                         -- read
			cpu_0_debug_mem_slave_readdata                      : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			cpu_0_debug_mem_slave_writedata                     : out std_logic_vector(31 downto 0);                     -- writedata
			cpu_0_debug_mem_slave_byteenable                    : out std_logic_vector(3 downto 0);                      -- byteenable
			cpu_0_debug_mem_slave_waitrequest                   : in  std_logic                      := 'X';             -- waitrequest
			cpu_0_debug_mem_slave_debugaccess                   : out std_logic;                                         -- debugaccess
			cpu_1_debug_mem_slave_address                       : out std_logic_vector(8 downto 0);                      -- address
			cpu_1_debug_mem_slave_write                         : out std_logic;                                         -- write
			cpu_1_debug_mem_slave_read                          : out std_logic;                                         -- read
			cpu_1_debug_mem_slave_readdata                      : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			cpu_1_debug_mem_slave_writedata                     : out std_logic_vector(31 downto 0);                     -- writedata
			cpu_1_debug_mem_slave_byteenable                    : out std_logic_vector(3 downto 0);                      -- byteenable
			cpu_1_debug_mem_slave_waitrequest                   : in  std_logic                      := 'X';             -- waitrequest
			cpu_1_debug_mem_slave_debugaccess                   : out std_logic;                                         -- debugaccess
			cpu_2_debug_mem_slave_address                       : out std_logic_vector(8 downto 0);                      -- address
			cpu_2_debug_mem_slave_write                         : out std_logic;                                         -- write
			cpu_2_debug_mem_slave_read                          : out std_logic;                                         -- read
			cpu_2_debug_mem_slave_readdata                      : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			cpu_2_debug_mem_slave_writedata                     : out std_logic_vector(31 downto 0);                     -- writedata
			cpu_2_debug_mem_slave_byteenable                    : out std_logic_vector(3 downto 0);                      -- byteenable
			cpu_2_debug_mem_slave_waitrequest                   : in  std_logic                      := 'X';             -- waitrequest
			cpu_2_debug_mem_slave_debugaccess                   : out std_logic;                                         -- debugaccess
			i2c_scl_s1_address                                  : out std_logic_vector(1 downto 0);                      -- address
			i2c_scl_s1_write                                    : out std_logic;                                         -- write
			i2c_scl_s1_readdata                                 : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			i2c_scl_s1_writedata                                : out std_logic_vector(31 downto 0);                     -- writedata
			i2c_scl_s1_chipselect                               : out std_logic;                                         -- chipselect
			i2c_sda_s1_address                                  : out std_logic_vector(1 downto 0);                      -- address
			i2c_sda_s1_write                                    : out std_logic;                                         -- write
			i2c_sda_s1_readdata                                 : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			i2c_sda_s1_writedata                                : out std_logic_vector(31 downto 0);                     -- writedata
			i2c_sda_s1_chipselect                               : out std_logic;                                         -- chipselect
			jtag_uart_0_avalon_jtag_slave_address               : out std_logic_vector(0 downto 0);                      -- address
			jtag_uart_0_avalon_jtag_slave_write                 : out std_logic;                                         -- write
			jtag_uart_0_avalon_jtag_slave_read                  : out std_logic;                                         -- read
			jtag_uart_0_avalon_jtag_slave_readdata              : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata             : out std_logic_vector(31 downto 0);                     -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest           : in  std_logic                      := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect            : out std_logic;                                         -- chipselect
			jtag_uart_1_avalon_jtag_slave_address               : out std_logic_vector(0 downto 0);                      -- address
			jtag_uart_1_avalon_jtag_slave_write                 : out std_logic;                                         -- write
			jtag_uart_1_avalon_jtag_slave_read                  : out std_logic;                                         -- read
			jtag_uart_1_avalon_jtag_slave_readdata              : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			jtag_uart_1_avalon_jtag_slave_writedata             : out std_logic_vector(31 downto 0);                     -- writedata
			jtag_uart_1_avalon_jtag_slave_waitrequest           : in  std_logic                      := 'X';             -- waitrequest
			jtag_uart_1_avalon_jtag_slave_chipselect            : out std_logic;                                         -- chipselect
			jtag_uart_2_avalon_jtag_slave_address               : out std_logic_vector(0 downto 0);                      -- address
			jtag_uart_2_avalon_jtag_slave_write                 : out std_logic;                                         -- write
			jtag_uart_2_avalon_jtag_slave_read                  : out std_logic;                                         -- read
			jtag_uart_2_avalon_jtag_slave_readdata              : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			jtag_uart_2_avalon_jtag_slave_writedata             : out std_logic_vector(31 downto 0);                     -- writedata
			jtag_uart_2_avalon_jtag_slave_waitrequest           : in  std_logic                      := 'X';             -- waitrequest
			jtag_uart_2_avalon_jtag_slave_chipselect            : out std_logic;                                         -- chipselect
			key_s1_address                                      : out std_logic_vector(1 downto 0);                      -- address
			key_s1_write                                        : out std_logic;                                         -- write
			key_s1_readdata                                     : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			key_s1_writedata                                    : out std_logic_vector(31 downto 0);                     -- writedata
			key_s1_chipselect                                   : out std_logic;                                         -- chipselect
			ledg_s1_address                                     : out std_logic_vector(2 downto 0);                      -- address
			ledg_s1_write                                       : out std_logic;                                         -- write
			ledg_s1_readdata                                    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			ledg_s1_writedata                                   : out std_logic_vector(31 downto 0);                     -- writedata
			ledg_s1_chipselect                                  : out std_logic;                                         -- chipselect
			ledr_s1_address                                     : out std_logic_vector(2 downto 0);                      -- address
			ledr_s1_write                                       : out std_logic;                                         -- write
			ledr_s1_readdata                                    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			ledr_s1_writedata                                   : out std_logic_vector(31 downto 0);                     -- writedata
			ledr_s1_chipselect                                  : out std_logic;                                         -- chipselect
			lpddr2_avl_0_address                                : out std_logic_vector(26 downto 0);                     -- address
			lpddr2_avl_0_write                                  : out std_logic;                                         -- write
			lpddr2_avl_0_read                                   : out std_logic;                                         -- read
			lpddr2_avl_0_readdata                               : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			lpddr2_avl_0_writedata                              : out std_logic_vector(31 downto 0);                     -- writedata
			lpddr2_avl_0_beginbursttransfer                     : out std_logic;                                         -- beginbursttransfer
			lpddr2_avl_0_burstcount                             : out std_logic_vector(7 downto 0);                      -- burstcount
			lpddr2_avl_0_byteenable                             : out std_logic_vector(3 downto 0);                      -- byteenable
			lpddr2_avl_0_readdatavalid                          : in  std_logic                      := 'X';             -- readdatavalid
			lpddr2_avl_0_waitrequest                            : in  std_logic                      := 'X';             -- waitrequest
			mailbox_simple_0_avmm_msg_receiver_address          : out std_logic_vector(1 downto 0);                      -- address
			mailbox_simple_0_avmm_msg_receiver_write            : out std_logic;                                         -- write
			mailbox_simple_0_avmm_msg_receiver_read             : out std_logic;                                         -- read
			mailbox_simple_0_avmm_msg_receiver_readdata         : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			mailbox_simple_0_avmm_msg_receiver_writedata        : out std_logic_vector(31 downto 0);                     -- writedata
			mailbox_simple_0_avmm_msg_sender_address            : out std_logic_vector(1 downto 0);                      -- address
			mailbox_simple_0_avmm_msg_sender_write              : out std_logic;                                         -- write
			mailbox_simple_0_avmm_msg_sender_read               : out std_logic;                                         -- read
			mailbox_simple_0_avmm_msg_sender_readdata           : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			mailbox_simple_0_avmm_msg_sender_writedata          : out std_logic_vector(31 downto 0);                     -- writedata
			mailbox_simple_0_avmm_msg_sender_waitrequest        : in  std_logic                      := 'X';             -- waitrequest
			mailbox_simple_1_avmm_msg_receiver_address          : out std_logic_vector(1 downto 0);                      -- address
			mailbox_simple_1_avmm_msg_receiver_write            : out std_logic;                                         -- write
			mailbox_simple_1_avmm_msg_receiver_read             : out std_logic;                                         -- read
			mailbox_simple_1_avmm_msg_receiver_readdata         : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			mailbox_simple_1_avmm_msg_receiver_writedata        : out std_logic_vector(31 downto 0);                     -- writedata
			mailbox_simple_1_avmm_msg_sender_address            : out std_logic_vector(1 downto 0);                      -- address
			mailbox_simple_1_avmm_msg_sender_write              : out std_logic;                                         -- write
			mailbox_simple_1_avmm_msg_sender_read               : out std_logic;                                         -- read
			mailbox_simple_1_avmm_msg_sender_readdata           : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			mailbox_simple_1_avmm_msg_sender_writedata          : out std_logic_vector(31 downto 0);                     -- writedata
			mailbox_simple_1_avmm_msg_sender_waitrequest        : in  std_logic                      := 'X';             -- waitrequest
			mailbox_simple_2_avmm_msg_receiver_address          : out std_logic_vector(1 downto 0);                      -- address
			mailbox_simple_2_avmm_msg_receiver_write            : out std_logic;                                         -- write
			mailbox_simple_2_avmm_msg_receiver_read             : out std_logic;                                         -- read
			mailbox_simple_2_avmm_msg_receiver_readdata         : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			mailbox_simple_2_avmm_msg_receiver_writedata        : out std_logic_vector(31 downto 0);                     -- writedata
			mailbox_simple_2_avmm_msg_sender_address            : out std_logic_vector(1 downto 0);                      -- address
			mailbox_simple_2_avmm_msg_sender_write              : out std_logic;                                         -- write
			mailbox_simple_2_avmm_msg_sender_read               : out std_logic;                                         -- read
			mailbox_simple_2_avmm_msg_sender_readdata           : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			mailbox_simple_2_avmm_msg_sender_writedata          : out std_logic_vector(31 downto 0);                     -- writedata
			mailbox_simple_2_avmm_msg_sender_waitrequest        : in  std_logic                      := 'X';             -- waitrequest
			mailbox_simple_3_avmm_msg_receiver_address          : out std_logic_vector(1 downto 0);                      -- address
			mailbox_simple_3_avmm_msg_receiver_write            : out std_logic;                                         -- write
			mailbox_simple_3_avmm_msg_receiver_read             : out std_logic;                                         -- read
			mailbox_simple_3_avmm_msg_receiver_readdata         : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			mailbox_simple_3_avmm_msg_receiver_writedata        : out std_logic_vector(31 downto 0);                     -- writedata
			mailbox_simple_3_avmm_msg_sender_address            : out std_logic_vector(1 downto 0);                      -- address
			mailbox_simple_3_avmm_msg_sender_write              : out std_logic;                                         -- write
			mailbox_simple_3_avmm_msg_sender_read               : out std_logic;                                         -- read
			mailbox_simple_3_avmm_msg_sender_readdata           : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			mailbox_simple_3_avmm_msg_sender_writedata          : out std_logic_vector(31 downto 0);                     -- writedata
			mailbox_simple_3_avmm_msg_sender_waitrequest        : in  std_logic                      := 'X';             -- waitrequest
			read_dma_0_csr_address                              : out std_logic_vector(2 downto 0);                      -- address
			read_dma_0_csr_write                                : out std_logic;                                         -- write
			read_dma_0_csr_read                                 : out std_logic;                                         -- read
			read_dma_0_csr_readdata                             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			read_dma_0_csr_writedata                            : out std_logic_vector(31 downto 0);                     -- writedata
			read_dma_0_csr_byteenable                           : out std_logic_vector(3 downto 0);                      -- byteenable
			read_dma_0_descriptor_slave_write                   : out std_logic;                                         -- write
			read_dma_0_descriptor_slave_writedata               : out std_logic_vector(127 downto 0);                    -- writedata
			read_dma_0_descriptor_slave_byteenable              : out std_logic_vector(15 downto 0);                     -- byteenable
			read_dma_0_descriptor_slave_waitrequest             : in  std_logic                      := 'X';             -- waitrequest
			sd_cont_0_slave_address                             : out std_logic_vector(7 downto 0);                      -- address
			sd_cont_0_slave_write                               : out std_logic;                                         -- write
			sd_cont_0_slave_read                                : out std_logic;                                         -- read
			sd_cont_0_slave_readdata                            : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			sd_cont_0_slave_writedata                           : out std_logic_vector(31 downto 0);                     -- writedata
			sd_cont_0_slave_waitrequest                         : in  std_logic                      := 'X';             -- waitrequest
			sd_cont_0_slave_chipselect                          : out std_logic;                                         -- chipselect
			sram_uas_address                                    : out std_logic_vector(18 downto 0);                     -- address
			sram_uas_write                                      : out std_logic;                                         -- write
			sram_uas_read                                       : out std_logic;                                         -- read
			sram_uas_readdata                                   : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- readdata
			sram_uas_writedata                                  : out std_logic_vector(15 downto 0);                     -- writedata
			sram_uas_burstcount                                 : out std_logic_vector(1 downto 0);                      -- burstcount
			sram_uas_byteenable                                 : out std_logic_vector(1 downto 0);                      -- byteenable
			sram_uas_readdatavalid                              : in  std_logic                      := 'X';             -- readdatavalid
			sram_uas_waitrequest                                : in  std_logic                      := 'X';             -- waitrequest
			sram_uas_lock                                       : out std_logic;                                         -- lock
			sram_uas_debugaccess                                : out std_logic;                                         -- debugaccess
			sysid_control_slave_address                         : out std_logic_vector(0 downto 0);                      -- address
			sysid_control_slave_readdata                        : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			timer_0_s1_address                                  : out std_logic_vector(2 downto 0);                      -- address
			timer_0_s1_write                                    : out std_logic;                                         -- write
			timer_0_s1_readdata                                 : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- readdata
			timer_0_s1_writedata                                : out std_logic_vector(15 downto 0);                     -- writedata
			timer_0_s1_chipselect                               : out std_logic;                                         -- chipselect
			timer_1_s1_address                                  : out std_logic_vector(3 downto 0);                      -- address
			timer_1_s1_write                                    : out std_logic;                                         -- write
			timer_1_s1_readdata                                 : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- readdata
			timer_1_s1_writedata                                : out std_logic_vector(15 downto 0);                     -- writedata
			timer_1_s1_chipselect                               : out std_logic;                                         -- chipselect
			video_dma_csr_address                               : out std_logic_vector(2 downto 0);                      -- address
			video_dma_csr_write                                 : out std_logic;                                         -- write
			video_dma_csr_read                                  : out std_logic;                                         -- read
			video_dma_csr_readdata                              : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			video_dma_csr_writedata                             : out std_logic_vector(31 downto 0);                     -- writedata
			video_dma_csr_byteenable                            : out std_logic_vector(3 downto 0);                      -- byteenable
			video_dma_descriptor_slave_write                    : out std_logic;                                         -- write
			video_dma_descriptor_slave_writedata                : out std_logic_vector(127 downto 0);                    -- writedata
			video_dma_descriptor_slave_byteenable               : out std_logic_vector(15 downto 0);                     -- byteenable
			video_dma_descriptor_slave_waitrequest              : in  std_logic                      := 'X';             -- waitrequest
			write_dma_0_csr_address                             : out std_logic_vector(2 downto 0);                      -- address
			write_dma_0_csr_write                               : out std_logic;                                         -- write
			write_dma_0_csr_read                                : out std_logic;                                         -- read
			write_dma_0_csr_readdata                            : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			write_dma_0_csr_writedata                           : out std_logic_vector(31 downto 0);                     -- writedata
			write_dma_0_csr_byteenable                          : out std_logic_vector(3 downto 0);                      -- byteenable
			write_dma_0_descriptor_slave_write                  : out std_logic;                                         -- write
			write_dma_0_descriptor_slave_writedata              : out std_logic_vector(127 downto 0);                    -- writedata
			write_dma_0_descriptor_slave_byteenable             : out std_logic_vector(15 downto 0);                     -- byteenable
			write_dma_0_descriptor_slave_waitrequest            : in  std_logic                      := 'X'              -- waitrequest
		);
	end component HW_QSYS_mm_interconnect_0;

	component HW_QSYS_mm_interconnect_1 is
		port (
			clk_125_clk_clk                                     : in  std_logic                     := 'X';             -- clk
			lpddr2_mp_cmd_reset_n_1_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			video_dma_reset_n_reset_bridge_in_reset_reset       : in  std_logic                     := 'X';             -- reset
			read_dma_0_mm_read_address                          : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			read_dma_0_mm_read_waitrequest                      : out std_logic;                                        -- waitrequest
			read_dma_0_mm_read_burstcount                       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- burstcount
			read_dma_0_mm_read_byteenable                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			read_dma_0_mm_read_read                             : in  std_logic                     := 'X';             -- read
			read_dma_0_mm_read_readdata                         : out std_logic_vector(31 downto 0);                    -- readdata
			read_dma_0_mm_read_readdatavalid                    : out std_logic;                                        -- readdatavalid
			video_dma_mm_read_address                           : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			video_dma_mm_read_waitrequest                       : out std_logic;                                        -- waitrequest
			video_dma_mm_read_burstcount                        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- burstcount
			video_dma_mm_read_byteenable                        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			video_dma_mm_read_read                              : in  std_logic                     := 'X';             -- read
			video_dma_mm_read_readdata                          : out std_logic_vector(31 downto 0);                    -- readdata
			video_dma_mm_read_readdatavalid                     : out std_logic;                                        -- readdatavalid
			lpddr2_avl_1_address                                : out std_logic_vector(26 downto 0);                    -- address
			lpddr2_avl_1_write                                  : out std_logic;                                        -- write
			lpddr2_avl_1_read                                   : out std_logic;                                        -- read
			lpddr2_avl_1_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			lpddr2_avl_1_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			lpddr2_avl_1_beginbursttransfer                     : out std_logic;                                        -- beginbursttransfer
			lpddr2_avl_1_burstcount                             : out std_logic_vector(7 downto 0);                     -- burstcount
			lpddr2_avl_1_byteenable                             : out std_logic_vector(3 downto 0);                     -- byteenable
			lpddr2_avl_1_readdatavalid                          : in  std_logic                     := 'X';             -- readdatavalid
			lpddr2_avl_1_waitrequest                            : in  std_logic                     := 'X'              -- waitrequest
		);
	end component HW_QSYS_mm_interconnect_1;

	component HW_QSYS_mm_interconnect_2 is
		port (
			clk_125_clk_clk                                     : in  std_logic                     := 'X';             -- clk
			lpddr2_mp_cmd_reset_n_2_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			write_dma_0_reset_n_reset_bridge_in_reset_reset     : in  std_logic                     := 'X';             -- reset
			write_dma_0_mm_write_address                        : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			write_dma_0_mm_write_waitrequest                    : out std_logic;                                        -- waitrequest
			write_dma_0_mm_write_burstcount                     : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- burstcount
			write_dma_0_mm_write_byteenable                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			write_dma_0_mm_write_write                          : in  std_logic                     := 'X';             -- write
			write_dma_0_mm_write_writedata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			lpddr2_avl_2_address                                : out std_logic_vector(26 downto 0);                    -- address
			lpddr2_avl_2_write                                  : out std_logic;                                        -- write
			lpddr2_avl_2_read                                   : out std_logic;                                        -- read
			lpddr2_avl_2_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			lpddr2_avl_2_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			lpddr2_avl_2_beginbursttransfer                     : out std_logic;                                        -- beginbursttransfer
			lpddr2_avl_2_burstcount                             : out std_logic_vector(7 downto 0);                     -- burstcount
			lpddr2_avl_2_byteenable                             : out std_logic_vector(3 downto 0);                     -- byteenable
			lpddr2_avl_2_readdatavalid                          : in  std_logic                     := 'X';             -- readdatavalid
			lpddr2_avl_2_waitrequest                            : in  std_logic                     := 'X'              -- waitrequest
		);
	end component HW_QSYS_mm_interconnect_2;

	component HW_QSYS_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			receiver5_irq : in  std_logic                     := 'X'; -- irq
			receiver6_irq : in  std_logic                     := 'X'; -- irq
			receiver7_irq : in  std_logic                     := 'X'; -- irq
			receiver8_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component HW_QSYS_irq_mapper;

	component HW_QSYS_irq_mapper_001 is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component HW_QSYS_irq_mapper_001;

	component HW_QSYS_avalon_st_adapter is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk        : in  std_logic                     := 'X';             -- clk
			in_rst_0_reset      : in  std_logic                     := 'X';             -- reset
			in_0_data           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_0_valid          : in  std_logic                     := 'X';             -- valid
			in_0_ready          : out std_logic;                                        -- ready
			in_0_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_0_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			in_0_empty          : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			out_0_data          : out std_logic_vector(31 downto 0);                    -- data
			out_0_valid         : out std_logic;                                        -- valid
			out_0_ready         : in  std_logic                     := 'X';             -- ready
			out_0_startofpacket : out std_logic;                                        -- startofpacket
			out_0_endofpacket   : out std_logic;                                        -- endofpacket
			out_0_empty         : out std_logic_vector(1 downto 0)                      -- empty
		);
	end component HW_QSYS_avalon_st_adapter;

	component HW_QSYS_avalon_st_adapter_001 is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk        : in  std_logic                     := 'X';             -- clk
			in_rst_0_reset      : in  std_logic                     := 'X';             -- reset
			in_0_data           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_0_valid          : in  std_logic                     := 'X';             -- valid
			in_0_ready          : out std_logic;                                        -- ready
			in_0_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_0_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			in_0_empty          : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			out_0_data          : out std_logic_vector(31 downto 0);                    -- data
			out_0_valid         : out std_logic;                                        -- valid
			out_0_ready         : in  std_logic                     := 'X';             -- ready
			out_0_startofpacket : out std_logic;                                        -- startofpacket
			out_0_endofpacket   : out std_logic;                                        -- endofpacket
			out_0_empty         : out std_logic_vector(1 downto 0)                      -- empty
		);
	end component HW_QSYS_avalon_st_adapter_001;

	component HW_qsys_reset_controller_0 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component HW_qsys_reset_controller_0;

	component HW_qsys_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component HW_qsys_rst_controller_001;

	signal twod_idct_st_hw_0_dst_valid                                     : std_logic;                      -- twod_idct_st_hw_0:dst_valid -> write_dma_0:st_sink_valid
	signal twod_idct_st_hw_0_dst_data                                      : std_logic_vector(31 downto 0);  -- twod_idct_st_hw_0:DATAOUT -> write_dma_0:st_sink_data
	signal twod_idct_st_hw_0_dst_ready                                     : std_logic;                      -- write_dma_0:st_sink_ready -> twod_idct_st_hw_0:dst_ready
	signal pixel_con_out_valid                                             : std_logic;                      -- Pixel_Con:valid_out -> video:valid
	signal pixel_con_out_data                                              : std_logic_vector(23 downto 0);  -- Pixel_Con:data_out -> video:data
	signal pixel_con_out_ready                                             : std_logic;                      -- video:ready -> Pixel_Con:ready_in
	signal pixel_con_out_startofpacket                                     : std_logic;                      -- Pixel_Con:sop_out -> video:sop
	signal pixel_con_out_endofpacket                                       : std_logic;                      -- Pixel_Con:eop_out -> video:eop
	signal pixel_con_out_empty                                             : std_logic;                      -- Pixel_Con:empty_out -> video:empty
	signal read_dma_0_st_source_valid                                      : std_logic;                      -- read_dma_0:st_source_valid -> twod_idct_st_hw_0:src_valid
	signal read_dma_0_st_source_data                                       : std_logic_vector(31 downto 0);  -- read_dma_0:st_source_data -> twod_idct_st_hw_0:DATAIN
	signal read_dma_0_st_source_ready                                      : std_logic;                      -- twod_idct_st_hw_0:src_ready -> read_dma_0:st_source_ready
	signal video_pll_outclk0_clk                                           : std_logic;                      -- video_pll:outclk_0 -> [video_clk_clk, Pixel_Con:clk, avalon_st_adapter:in_clk_0_clk, rst_controller:clk, video:clk, video_fifo:rdclock]
	signal reset_controller_0_reset_out_reset                              : std_logic;                      -- reset_controller_0:reset_out -> [reset_controller_0_reset_out_reset:in, rst_controller:reset_in0, rst_controller_001:reset_in1, rst_controller_002:reset_in1, rst_controller_003:reset_in1, rst_controller_004:reset_in0, rst_controller_005:reset_in0, video_pll:rst]
	signal sram_sharer_tcm_request                                         : std_logic;                      -- sram_sharer:request -> sram_bridge:request
	signal sram_sharer_tcm_sram_tcm_byteenable_n_out_out                   : std_logic_vector(1 downto 0);   -- sram_sharer:sram_tcm_byteenable_n_out -> sram_bridge:tcs_sram_tcm_byteenable_n_out
	signal sram_sharer_tcm_sram_tcm_data_out_outen                         : std_logic;                      -- sram_sharer:sram_tcm_data_outen -> sram_bridge:tcs_sram_tcm_data_outen
	signal sram_sharer_tcm_sram_tcm_data_out_in                            : std_logic_vector(15 downto 0);  -- sram_bridge:tcs_sram_tcm_data_in -> sram_sharer:sram_tcm_data_in
	signal sram_sharer_tcm_sram_tcm_write_n_out_out                        : std_logic_vector(0 downto 0);   -- sram_sharer:sram_tcm_write_n_out -> sram_bridge:tcs_sram_tcm_write_n_out
	signal sram_sharer_tcm_sram_tcm_data_out_out                           : std_logic_vector(15 downto 0);  -- sram_sharer:sram_tcm_data_out -> sram_bridge:tcs_sram_tcm_data_out
	signal sram_sharer_tcm_sram_tcm_address_out_out                        : std_logic_vector(18 downto 0);  -- sram_sharer:sram_tcm_address_out -> sram_bridge:tcs_sram_tcm_address_out
	signal sram_sharer_tcm_sram_tcm_chipselect_n_out_out                   : std_logic_vector(0 downto 0);   -- sram_sharer:sram_tcm_chipselect_n_out -> sram_bridge:tcs_sram_tcm_chipselect_n_out
	signal sram_sharer_tcm_grant                                           : std_logic;                      -- sram_bridge:grant -> sram_sharer:grant
	signal sram_sharer_tcm_sram_tcm_outputenable_n_out_out                 : std_logic_vector(0 downto 0);   -- sram_sharer:sram_tcm_outputenable_n_out -> sram_bridge:tcs_sram_tcm_outputenable_n_out
	signal sram_tcm_data_outen                                             : std_logic;                      -- sram:tcm_data_outen -> sram_sharer:tcs0_data_outen
	signal sram_tcm_outputenable_n_out                                     : std_logic;                      -- sram:tcm_outputenable_n_out -> sram_sharer:tcs0_outputenable_n_out
	signal sram_tcm_request                                                : std_logic;                      -- sram:tcm_request -> sram_sharer:tcs0_request
	signal sram_tcm_byteenable_n_out                                       : std_logic_vector(1 downto 0);   -- sram:tcm_byteenable_n_out -> sram_sharer:tcs0_byteenable_n_out
	signal sram_tcm_write_n_out                                            : std_logic;                      -- sram:tcm_write_n_out -> sram_sharer:tcs0_write_n_out
	signal sram_tcm_grant                                                  : std_logic;                      -- sram_sharer:tcs0_grant -> sram:tcm_grant
	signal sram_tcm_chipselect_n_out                                       : std_logic;                      -- sram:tcm_chipselect_n_out -> sram_sharer:tcs0_chipselect_n_out
	signal sram_tcm_address_out                                            : std_logic_vector(18 downto 0);  -- sram:tcm_address_out -> sram_sharer:tcs0_address_out
	signal sram_tcm_data_out                                               : std_logic_vector(15 downto 0);  -- sram:tcm_data_out -> sram_sharer:tcs0_data_out
	signal sram_tcm_data_in                                                : std_logic_vector(15 downto 0);  -- sram_sharer:tcs0_data_in -> sram:tcm_data_in
	signal cpu_0_data_master_readdata                                      : std_logic_vector(31 downto 0);  -- mm_interconnect_0:cpu_0_data_master_readdata -> cpu_0:d_readdata
	signal cpu_0_data_master_waitrequest                                   : std_logic;                      -- mm_interconnect_0:cpu_0_data_master_waitrequest -> cpu_0:d_waitrequest
	signal cpu_0_data_master_debugaccess                                   : std_logic;                      -- cpu_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_0_data_master_debugaccess
	signal cpu_0_data_master_address                                       : std_logic_vector(29 downto 0);  -- cpu_0:d_address -> mm_interconnect_0:cpu_0_data_master_address
	signal cpu_0_data_master_byteenable                                    : std_logic_vector(3 downto 0);   -- cpu_0:d_byteenable -> mm_interconnect_0:cpu_0_data_master_byteenable
	signal cpu_0_data_master_read                                          : std_logic;                      -- cpu_0:d_read -> mm_interconnect_0:cpu_0_data_master_read
	signal cpu_0_data_master_readdatavalid                                 : std_logic;                      -- mm_interconnect_0:cpu_0_data_master_readdatavalid -> cpu_0:d_readdatavalid
	signal cpu_0_data_master_write                                         : std_logic;                      -- cpu_0:d_write -> mm_interconnect_0:cpu_0_data_master_write
	signal cpu_0_data_master_writedata                                     : std_logic_vector(31 downto 0);  -- cpu_0:d_writedata -> mm_interconnect_0:cpu_0_data_master_writedata
	signal cpu_0_data_master_burstcount                                    : std_logic_vector(3 downto 0);   -- cpu_0:d_burstcount -> mm_interconnect_0:cpu_0_data_master_burstcount
	signal cpu_1_data_master_readdata                                      : std_logic_vector(31 downto 0);  -- mm_interconnect_0:cpu_1_data_master_readdata -> cpu_1:d_readdata
	signal cpu_1_data_master_waitrequest                                   : std_logic;                      -- mm_interconnect_0:cpu_1_data_master_waitrequest -> cpu_1:d_waitrequest
	signal cpu_1_data_master_debugaccess                                   : std_logic;                      -- cpu_1:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_1_data_master_debugaccess
	signal cpu_1_data_master_address                                       : std_logic_vector(29 downto 0);  -- cpu_1:d_address -> mm_interconnect_0:cpu_1_data_master_address
	signal cpu_1_data_master_byteenable                                    : std_logic_vector(3 downto 0);   -- cpu_1:d_byteenable -> mm_interconnect_0:cpu_1_data_master_byteenable
	signal cpu_1_data_master_read                                          : std_logic;                      -- cpu_1:d_read -> mm_interconnect_0:cpu_1_data_master_read
	signal cpu_1_data_master_readdatavalid                                 : std_logic;                      -- mm_interconnect_0:cpu_1_data_master_readdatavalid -> cpu_1:d_readdatavalid
	signal cpu_1_data_master_write                                         : std_logic;                      -- cpu_1:d_write -> mm_interconnect_0:cpu_1_data_master_write
	signal cpu_1_data_master_writedata                                     : std_logic_vector(31 downto 0);  -- cpu_1:d_writedata -> mm_interconnect_0:cpu_1_data_master_writedata
	signal cpu_1_data_master_burstcount                                    : std_logic_vector(3 downto 0);   -- cpu_1:d_burstcount -> mm_interconnect_0:cpu_1_data_master_burstcount
	signal cpu_2_data_master_readdata                                      : std_logic_vector(31 downto 0);  -- mm_interconnect_0:cpu_2_data_master_readdata -> cpu_2:d_readdata
	signal cpu_2_data_master_waitrequest                                   : std_logic;                      -- mm_interconnect_0:cpu_2_data_master_waitrequest -> cpu_2:d_waitrequest
	signal cpu_2_data_master_debugaccess                                   : std_logic;                      -- cpu_2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_2_data_master_debugaccess
	signal cpu_2_data_master_address                                       : std_logic_vector(29 downto 0);  -- cpu_2:d_address -> mm_interconnect_0:cpu_2_data_master_address
	signal cpu_2_data_master_byteenable                                    : std_logic_vector(3 downto 0);   -- cpu_2:d_byteenable -> mm_interconnect_0:cpu_2_data_master_byteenable
	signal cpu_2_data_master_read                                          : std_logic;                      -- cpu_2:d_read -> mm_interconnect_0:cpu_2_data_master_read
	signal cpu_2_data_master_readdatavalid                                 : std_logic;                      -- mm_interconnect_0:cpu_2_data_master_readdatavalid -> cpu_2:d_readdatavalid
	signal cpu_2_data_master_write                                         : std_logic;                      -- cpu_2:d_write -> mm_interconnect_0:cpu_2_data_master_write
	signal cpu_2_data_master_writedata                                     : std_logic_vector(31 downto 0);  -- cpu_2:d_writedata -> mm_interconnect_0:cpu_2_data_master_writedata
	signal cpu_2_data_master_burstcount                                    : std_logic_vector(3 downto 0);   -- cpu_2:d_burstcount -> mm_interconnect_0:cpu_2_data_master_burstcount
	signal cpu_0_instruction_master_readdata                               : std_logic_vector(31 downto 0);  -- mm_interconnect_0:cpu_0_instruction_master_readdata -> cpu_0:i_readdata
	signal cpu_0_instruction_master_waitrequest                            : std_logic;                      -- mm_interconnect_0:cpu_0_instruction_master_waitrequest -> cpu_0:i_waitrequest
	signal cpu_0_instruction_master_address                                : std_logic_vector(29 downto 0);  -- cpu_0:i_address -> mm_interconnect_0:cpu_0_instruction_master_address
	signal cpu_0_instruction_master_read                                   : std_logic;                      -- cpu_0:i_read -> mm_interconnect_0:cpu_0_instruction_master_read
	signal cpu_0_instruction_master_readdatavalid                          : std_logic;                      -- mm_interconnect_0:cpu_0_instruction_master_readdatavalid -> cpu_0:i_readdatavalid
	signal cpu_1_instruction_master_readdata                               : std_logic_vector(31 downto 0);  -- mm_interconnect_0:cpu_1_instruction_master_readdata -> cpu_1:i_readdata
	signal cpu_1_instruction_master_waitrequest                            : std_logic;                      -- mm_interconnect_0:cpu_1_instruction_master_waitrequest -> cpu_1:i_waitrequest
	signal cpu_1_instruction_master_address                                : std_logic_vector(29 downto 0);  -- cpu_1:i_address -> mm_interconnect_0:cpu_1_instruction_master_address
	signal cpu_1_instruction_master_read                                   : std_logic;                      -- cpu_1:i_read -> mm_interconnect_0:cpu_1_instruction_master_read
	signal cpu_1_instruction_master_readdatavalid                          : std_logic;                      -- mm_interconnect_0:cpu_1_instruction_master_readdatavalid -> cpu_1:i_readdatavalid
	signal cpu_2_instruction_master_readdata                               : std_logic_vector(31 downto 0);  -- mm_interconnect_0:cpu_2_instruction_master_readdata -> cpu_2:i_readdata
	signal cpu_2_instruction_master_waitrequest                            : std_logic;                      -- mm_interconnect_0:cpu_2_instruction_master_waitrequest -> cpu_2:i_waitrequest
	signal cpu_2_instruction_master_address                                : std_logic_vector(29 downto 0);  -- cpu_2:i_address -> mm_interconnect_0:cpu_2_instruction_master_address
	signal cpu_2_instruction_master_read                                   : std_logic;                      -- cpu_2:i_read -> mm_interconnect_0:cpu_2_instruction_master_read
	signal cpu_2_instruction_master_readdatavalid                          : std_logic;                      -- mm_interconnect_0:cpu_2_instruction_master_readdatavalid -> cpu_2:i_readdatavalid
	signal sd_cont_0_master_readdata                                       : std_logic_vector(31 downto 0);  -- mm_interconnect_0:sd_cont_0_master_readdata -> sd_cont_0:m_readdata
	signal mm_interconnect_0_sd_cont_0_master_waitrequest                  : std_logic;                      -- mm_interconnect_0:sd_cont_0_master_waitrequest -> mm_interconnect_0_sd_cont_0_master_waitrequest:in
	signal sd_cont_0_master_address                                        : std_logic_vector(31 downto 0);  -- sd_cont_0:m_address -> mm_interconnect_0:sd_cont_0_master_address
	signal sd_cont_0_master_read                                           : std_logic;                      -- sd_cont_0:m_read -> mm_interconnect_0:sd_cont_0_master_read
	signal sd_cont_0_master_write                                          : std_logic;                      -- sd_cont_0:m_write -> mm_interconnect_0:sd_cont_0_master_write
	signal sd_cont_0_master_writedata                                      : std_logic_vector(31 downto 0);  -- sd_cont_0:m_writedata -> mm_interconnect_0:sd_cont_0_master_writedata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect      : std_logic;                      -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0);  -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest     : std_logic;                      -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);   -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read            : std_logic;                      -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write           : std_logic;                      -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_lpddr2_avl_0_beginbursttransfer               : std_logic;                      -- mm_interconnect_0:lpddr2_avl_0_beginbursttransfer -> lpddr2:avl_burstbegin_0
	signal mm_interconnect_0_lpddr2_avl_0_readdata                         : std_logic_vector(31 downto 0);  -- lpddr2:avl_rdata_0 -> mm_interconnect_0:lpddr2_avl_0_readdata
	signal lpddr2_avl_0_waitrequest                                        : std_logic;                      -- lpddr2:avl_ready_0 -> lpddr2_avl_0_waitrequest:in
	signal mm_interconnect_0_lpddr2_avl_0_address                          : std_logic_vector(26 downto 0);  -- mm_interconnect_0:lpddr2_avl_0_address -> lpddr2:avl_addr_0
	signal mm_interconnect_0_lpddr2_avl_0_read                             : std_logic;                      -- mm_interconnect_0:lpddr2_avl_0_read -> lpddr2:avl_read_req_0
	signal mm_interconnect_0_lpddr2_avl_0_byteenable                       : std_logic_vector(3 downto 0);   -- mm_interconnect_0:lpddr2_avl_0_byteenable -> lpddr2:avl_be_0
	signal mm_interconnect_0_lpddr2_avl_0_readdatavalid                    : std_logic;                      -- lpddr2:avl_rdata_valid_0 -> mm_interconnect_0:lpddr2_avl_0_readdatavalid
	signal mm_interconnect_0_lpddr2_avl_0_write                            : std_logic;                      -- mm_interconnect_0:lpddr2_avl_0_write -> lpddr2:avl_write_req_0
	signal mm_interconnect_0_lpddr2_avl_0_writedata                        : std_logic_vector(31 downto 0);  -- mm_interconnect_0:lpddr2_avl_0_writedata -> lpddr2:avl_wdata_0
	signal mm_interconnect_0_lpddr2_avl_0_burstcount                       : std_logic_vector(7 downto 0);   -- mm_interconnect_0:lpddr2_avl_0_burstcount -> lpddr2:avl_size_0
	signal mm_interconnect_0_mailbox_simple_1_avmm_msg_receiver_readdata   : std_logic_vector(31 downto 0);  -- mailbox_simple_1:avmm_rcv_readdata -> mm_interconnect_0:mailbox_simple_1_avmm_msg_receiver_readdata
	signal mm_interconnect_0_mailbox_simple_1_avmm_msg_receiver_address    : std_logic_vector(1 downto 0);   -- mm_interconnect_0:mailbox_simple_1_avmm_msg_receiver_address -> mailbox_simple_1:avmm_rcv_address
	signal mm_interconnect_0_mailbox_simple_1_avmm_msg_receiver_read       : std_logic;                      -- mm_interconnect_0:mailbox_simple_1_avmm_msg_receiver_read -> mailbox_simple_1:avmm_rcv_read
	signal mm_interconnect_0_mailbox_simple_1_avmm_msg_receiver_write      : std_logic;                      -- mm_interconnect_0:mailbox_simple_1_avmm_msg_receiver_write -> mailbox_simple_1:avmm_rcv_write
	signal mm_interconnect_0_mailbox_simple_1_avmm_msg_receiver_writedata  : std_logic_vector(31 downto 0);  -- mm_interconnect_0:mailbox_simple_1_avmm_msg_receiver_writedata -> mailbox_simple_1:avmm_rcv_writedata
	signal mm_interconnect_0_mailbox_simple_2_avmm_msg_receiver_readdata   : std_logic_vector(31 downto 0);  -- mailbox_simple_2:avmm_rcv_readdata -> mm_interconnect_0:mailbox_simple_2_avmm_msg_receiver_readdata
	signal mm_interconnect_0_mailbox_simple_2_avmm_msg_receiver_address    : std_logic_vector(1 downto 0);   -- mm_interconnect_0:mailbox_simple_2_avmm_msg_receiver_address -> mailbox_simple_2:avmm_rcv_address
	signal mm_interconnect_0_mailbox_simple_2_avmm_msg_receiver_read       : std_logic;                      -- mm_interconnect_0:mailbox_simple_2_avmm_msg_receiver_read -> mailbox_simple_2:avmm_rcv_read
	signal mm_interconnect_0_mailbox_simple_2_avmm_msg_receiver_write      : std_logic;                      -- mm_interconnect_0:mailbox_simple_2_avmm_msg_receiver_write -> mailbox_simple_2:avmm_rcv_write
	signal mm_interconnect_0_mailbox_simple_2_avmm_msg_receiver_writedata  : std_logic_vector(31 downto 0);  -- mm_interconnect_0:mailbox_simple_2_avmm_msg_receiver_writedata -> mailbox_simple_2:avmm_rcv_writedata
	signal mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_readdata     : std_logic_vector(31 downto 0);  -- mailbox_simple_0:avmm_snd_readdata -> mm_interconnect_0:mailbox_simple_0_avmm_msg_sender_readdata
	signal mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_waitrequest  : std_logic;                      -- mailbox_simple_0:avmm_snd_waitrequest -> mm_interconnect_0:mailbox_simple_0_avmm_msg_sender_waitrequest
	signal mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_address      : std_logic_vector(1 downto 0);   -- mm_interconnect_0:mailbox_simple_0_avmm_msg_sender_address -> mailbox_simple_0:avmm_snd_address
	signal mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_read         : std_logic;                      -- mm_interconnect_0:mailbox_simple_0_avmm_msg_sender_read -> mailbox_simple_0:avmm_snd_read
	signal mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_write        : std_logic;                      -- mm_interconnect_0:mailbox_simple_0_avmm_msg_sender_write -> mailbox_simple_0:avmm_snd_write
	signal mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_writedata    : std_logic_vector(31 downto 0);  -- mm_interconnect_0:mailbox_simple_0_avmm_msg_sender_writedata -> mailbox_simple_0:avmm_snd_writedata
	signal mm_interconnect_0_mailbox_simple_3_avmm_msg_sender_readdata     : std_logic_vector(31 downto 0);  -- mailbox_simple_3:avmm_snd_readdata -> mm_interconnect_0:mailbox_simple_3_avmm_msg_sender_readdata
	signal mm_interconnect_0_mailbox_simple_3_avmm_msg_sender_waitrequest  : std_logic;                      -- mailbox_simple_3:avmm_snd_waitrequest -> mm_interconnect_0:mailbox_simple_3_avmm_msg_sender_waitrequest
	signal mm_interconnect_0_mailbox_simple_3_avmm_msg_sender_address      : std_logic_vector(1 downto 0);   -- mm_interconnect_0:mailbox_simple_3_avmm_msg_sender_address -> mailbox_simple_3:avmm_snd_address
	signal mm_interconnect_0_mailbox_simple_3_avmm_msg_sender_read         : std_logic;                      -- mm_interconnect_0:mailbox_simple_3_avmm_msg_sender_read -> mailbox_simple_3:avmm_snd_read
	signal mm_interconnect_0_mailbox_simple_3_avmm_msg_sender_write        : std_logic;                      -- mm_interconnect_0:mailbox_simple_3_avmm_msg_sender_write -> mailbox_simple_3:avmm_snd_write
	signal mm_interconnect_0_mailbox_simple_3_avmm_msg_sender_writedata    : std_logic_vector(31 downto 0);  -- mm_interconnect_0:mailbox_simple_3_avmm_msg_sender_writedata -> mailbox_simple_3:avmm_snd_writedata
	signal mm_interconnect_0_sysid_control_slave_readdata                  : std_logic_vector(31 downto 0);  -- sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	signal mm_interconnect_0_sysid_control_slave_address                   : std_logic_vector(0 downto 0);   -- mm_interconnect_0:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_0_video_dma_csr_readdata                        : std_logic_vector(31 downto 0);  -- video_dma:csr_readdata -> mm_interconnect_0:video_dma_csr_readdata
	signal mm_interconnect_0_video_dma_csr_address                         : std_logic_vector(2 downto 0);   -- mm_interconnect_0:video_dma_csr_address -> video_dma:csr_address
	signal mm_interconnect_0_video_dma_csr_read                            : std_logic;                      -- mm_interconnect_0:video_dma_csr_read -> video_dma:csr_read
	signal mm_interconnect_0_video_dma_csr_byteenable                      : std_logic_vector(3 downto 0);   -- mm_interconnect_0:video_dma_csr_byteenable -> video_dma:csr_byteenable
	signal mm_interconnect_0_video_dma_csr_write                           : std_logic;                      -- mm_interconnect_0:video_dma_csr_write -> video_dma:csr_write
	signal mm_interconnect_0_video_dma_csr_writedata                       : std_logic_vector(31 downto 0);  -- mm_interconnect_0:video_dma_csr_writedata -> video_dma:csr_writedata
	signal mm_interconnect_0_write_dma_0_csr_readdata                      : std_logic_vector(31 downto 0);  -- write_dma_0:csr_readdata -> mm_interconnect_0:write_dma_0_csr_readdata
	signal mm_interconnect_0_write_dma_0_csr_address                       : std_logic_vector(2 downto 0);   -- mm_interconnect_0:write_dma_0_csr_address -> write_dma_0:csr_address
	signal mm_interconnect_0_write_dma_0_csr_read                          : std_logic;                      -- mm_interconnect_0:write_dma_0_csr_read -> write_dma_0:csr_read
	signal mm_interconnect_0_write_dma_0_csr_byteenable                    : std_logic_vector(3 downto 0);   -- mm_interconnect_0:write_dma_0_csr_byteenable -> write_dma_0:csr_byteenable
	signal mm_interconnect_0_write_dma_0_csr_write                         : std_logic;                      -- mm_interconnect_0:write_dma_0_csr_write -> write_dma_0:csr_write
	signal mm_interconnect_0_write_dma_0_csr_writedata                     : std_logic_vector(31 downto 0);  -- mm_interconnect_0:write_dma_0_csr_writedata -> write_dma_0:csr_writedata
	signal mm_interconnect_0_read_dma_0_csr_readdata                       : std_logic_vector(31 downto 0);  -- read_dma_0:csr_readdata -> mm_interconnect_0:read_dma_0_csr_readdata
	signal mm_interconnect_0_read_dma_0_csr_address                        : std_logic_vector(2 downto 0);   -- mm_interconnect_0:read_dma_0_csr_address -> read_dma_0:csr_address
	signal mm_interconnect_0_read_dma_0_csr_read                           : std_logic;                      -- mm_interconnect_0:read_dma_0_csr_read -> read_dma_0:csr_read
	signal mm_interconnect_0_read_dma_0_csr_byteenable                     : std_logic_vector(3 downto 0);   -- mm_interconnect_0:read_dma_0_csr_byteenable -> read_dma_0:csr_byteenable
	signal mm_interconnect_0_read_dma_0_csr_write                          : std_logic;                      -- mm_interconnect_0:read_dma_0_csr_write -> read_dma_0:csr_write
	signal mm_interconnect_0_read_dma_0_csr_writedata                      : std_logic_vector(31 downto 0);  -- mm_interconnect_0:read_dma_0_csr_writedata -> read_dma_0:csr_writedata
	signal mm_interconnect_0_cpu_0_debug_mem_slave_readdata                : std_logic_vector(31 downto 0);  -- cpu_0:debug_mem_slave_readdata -> mm_interconnect_0:cpu_0_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest             : std_logic;                      -- cpu_0:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess             : std_logic;                      -- mm_interconnect_0:cpu_0_debug_mem_slave_debugaccess -> cpu_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_0_debug_mem_slave_address                 : std_logic_vector(8 downto 0);   -- mm_interconnect_0:cpu_0_debug_mem_slave_address -> cpu_0:debug_mem_slave_address
	signal mm_interconnect_0_cpu_0_debug_mem_slave_read                    : std_logic;                      -- mm_interconnect_0:cpu_0_debug_mem_slave_read -> cpu_0:debug_mem_slave_read
	signal mm_interconnect_0_cpu_0_debug_mem_slave_byteenable              : std_logic_vector(3 downto 0);   -- mm_interconnect_0:cpu_0_debug_mem_slave_byteenable -> cpu_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_0_debug_mem_slave_write                   : std_logic;                      -- mm_interconnect_0:cpu_0_debug_mem_slave_write -> cpu_0:debug_mem_slave_write
	signal mm_interconnect_0_cpu_0_debug_mem_slave_writedata               : std_logic_vector(31 downto 0);  -- mm_interconnect_0:cpu_0_debug_mem_slave_writedata -> cpu_0:debug_mem_slave_writedata
	signal mm_interconnect_0_video_dma_descriptor_slave_waitrequest        : std_logic;                      -- video_dma:descriptor_slave_waitrequest -> mm_interconnect_0:video_dma_descriptor_slave_waitrequest
	signal mm_interconnect_0_video_dma_descriptor_slave_byteenable         : std_logic_vector(15 downto 0);  -- mm_interconnect_0:video_dma_descriptor_slave_byteenable -> video_dma:descriptor_slave_byteenable
	signal mm_interconnect_0_video_dma_descriptor_slave_write              : std_logic;                      -- mm_interconnect_0:video_dma_descriptor_slave_write -> video_dma:descriptor_slave_write
	signal mm_interconnect_0_video_dma_descriptor_slave_writedata          : std_logic_vector(127 downto 0); -- mm_interconnect_0:video_dma_descriptor_slave_writedata -> video_dma:descriptor_slave_writedata
	signal mm_interconnect_0_write_dma_0_descriptor_slave_waitrequest      : std_logic;                      -- write_dma_0:descriptor_slave_waitrequest -> mm_interconnect_0:write_dma_0_descriptor_slave_waitrequest
	signal mm_interconnect_0_write_dma_0_descriptor_slave_byteenable       : std_logic_vector(15 downto 0);  -- mm_interconnect_0:write_dma_0_descriptor_slave_byteenable -> write_dma_0:descriptor_slave_byteenable
	signal mm_interconnect_0_write_dma_0_descriptor_slave_write            : std_logic;                      -- mm_interconnect_0:write_dma_0_descriptor_slave_write -> write_dma_0:descriptor_slave_write
	signal mm_interconnect_0_write_dma_0_descriptor_slave_writedata        : std_logic_vector(127 downto 0); -- mm_interconnect_0:write_dma_0_descriptor_slave_writedata -> write_dma_0:descriptor_slave_writedata
	signal mm_interconnect_0_read_dma_0_descriptor_slave_waitrequest       : std_logic;                      -- read_dma_0:descriptor_slave_waitrequest -> mm_interconnect_0:read_dma_0_descriptor_slave_waitrequest
	signal mm_interconnect_0_read_dma_0_descriptor_slave_byteenable        : std_logic_vector(15 downto 0);  -- mm_interconnect_0:read_dma_0_descriptor_slave_byteenable -> read_dma_0:descriptor_slave_byteenable
	signal mm_interconnect_0_read_dma_0_descriptor_slave_write             : std_logic;                      -- mm_interconnect_0:read_dma_0_descriptor_slave_write -> read_dma_0:descriptor_slave_write
	signal mm_interconnect_0_read_dma_0_descriptor_slave_writedata         : std_logic_vector(127 downto 0); -- mm_interconnect_0:read_dma_0_descriptor_slave_writedata -> read_dma_0:descriptor_slave_writedata
	signal mm_interconnect_0_timer_0_s1_chipselect                         : std_logic;                      -- mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	signal mm_interconnect_0_timer_0_s1_readdata                           : std_logic_vector(15 downto 0);  -- timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	signal mm_interconnect_0_timer_0_s1_address                            : std_logic_vector(2 downto 0);   -- mm_interconnect_0:timer_0_s1_address -> timer_0:address
	signal mm_interconnect_0_timer_0_s1_write                              : std_logic;                      -- mm_interconnect_0:timer_0_s1_write -> mm_interconnect_0_timer_0_s1_write:in
	signal mm_interconnect_0_timer_0_s1_writedata                          : std_logic_vector(15 downto 0);  -- mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	signal mm_interconnect_0_key_s1_chipselect                             : std_logic;                      -- mm_interconnect_0:key_s1_chipselect -> key:chipselect
	signal mm_interconnect_0_key_s1_readdata                               : std_logic_vector(31 downto 0);  -- key:readdata -> mm_interconnect_0:key_s1_readdata
	signal mm_interconnect_0_key_s1_address                                : std_logic_vector(1 downto 0);   -- mm_interconnect_0:key_s1_address -> key:address
	signal mm_interconnect_0_key_s1_write                                  : std_logic;                      -- mm_interconnect_0:key_s1_write -> mm_interconnect_0_key_s1_write:in
	signal mm_interconnect_0_key_s1_writedata                              : std_logic_vector(31 downto 0);  -- mm_interconnect_0:key_s1_writedata -> key:writedata
	signal mm_interconnect_0_timer_1_s1_chipselect                         : std_logic;                      -- mm_interconnect_0:timer_1_s1_chipselect -> timer_1:chipselect
	signal mm_interconnect_0_timer_1_s1_readdata                           : std_logic_vector(15 downto 0);  -- timer_1:readdata -> mm_interconnect_0:timer_1_s1_readdata
	signal mm_interconnect_0_timer_1_s1_address                            : std_logic_vector(3 downto 0);   -- mm_interconnect_0:timer_1_s1_address -> timer_1:address
	signal mm_interconnect_0_timer_1_s1_write                              : std_logic;                      -- mm_interconnect_0:timer_1_s1_write -> mm_interconnect_0_timer_1_s1_write:in
	signal mm_interconnect_0_timer_1_s1_writedata                          : std_logic_vector(15 downto 0);  -- mm_interconnect_0:timer_1_s1_writedata -> timer_1:writedata
	signal mm_interconnect_0_ledg_s1_chipselect                            : std_logic;                      -- mm_interconnect_0:ledg_s1_chipselect -> ledg:chipselect
	signal mm_interconnect_0_ledg_s1_readdata                              : std_logic_vector(31 downto 0);  -- ledg:readdata -> mm_interconnect_0:ledg_s1_readdata
	signal mm_interconnect_0_ledg_s1_address                               : std_logic_vector(2 downto 0);   -- mm_interconnect_0:ledg_s1_address -> ledg:address
	signal mm_interconnect_0_ledg_s1_write                                 : std_logic;                      -- mm_interconnect_0:ledg_s1_write -> mm_interconnect_0_ledg_s1_write:in
	signal mm_interconnect_0_ledg_s1_writedata                             : std_logic_vector(31 downto 0);  -- mm_interconnect_0:ledg_s1_writedata -> ledg:writedata
	signal mm_interconnect_0_ledr_s1_chipselect                            : std_logic;                      -- mm_interconnect_0:ledr_s1_chipselect -> ledr:chipselect
	signal mm_interconnect_0_ledr_s1_readdata                              : std_logic_vector(31 downto 0);  -- ledr:readdata -> mm_interconnect_0:ledr_s1_readdata
	signal mm_interconnect_0_ledr_s1_address                               : std_logic_vector(2 downto 0);   -- mm_interconnect_0:ledr_s1_address -> ledr:address
	signal mm_interconnect_0_ledr_s1_write                                 : std_logic;                      -- mm_interconnect_0:ledr_s1_write -> mm_interconnect_0_ledr_s1_write:in
	signal mm_interconnect_0_ledr_s1_writedata                             : std_logic_vector(31 downto 0);  -- mm_interconnect_0:ledr_s1_writedata -> ledr:writedata
	signal mm_interconnect_0_i2c_scl_s1_chipselect                         : std_logic;                      -- mm_interconnect_0:i2c_scl_s1_chipselect -> i2c_scl:chipselect
	signal mm_interconnect_0_i2c_scl_s1_readdata                           : std_logic_vector(31 downto 0);  -- i2c_scl:readdata -> mm_interconnect_0:i2c_scl_s1_readdata
	signal mm_interconnect_0_i2c_scl_s1_address                            : std_logic_vector(1 downto 0);   -- mm_interconnect_0:i2c_scl_s1_address -> i2c_scl:address
	signal mm_interconnect_0_i2c_scl_s1_write                              : std_logic;                      -- mm_interconnect_0:i2c_scl_s1_write -> mm_interconnect_0_i2c_scl_s1_write:in
	signal mm_interconnect_0_i2c_scl_s1_writedata                          : std_logic_vector(31 downto 0);  -- mm_interconnect_0:i2c_scl_s1_writedata -> i2c_scl:writedata
	signal mm_interconnect_0_i2c_sda_s1_chipselect                         : std_logic;                      -- mm_interconnect_0:i2c_sda_s1_chipselect -> i2c_sda:chipselect
	signal mm_interconnect_0_i2c_sda_s1_readdata                           : std_logic_vector(31 downto 0);  -- i2c_sda:readdata -> mm_interconnect_0:i2c_sda_s1_readdata
	signal mm_interconnect_0_i2c_sda_s1_address                            : std_logic_vector(1 downto 0);   -- mm_interconnect_0:i2c_sda_s1_address -> i2c_sda:address
	signal mm_interconnect_0_i2c_sda_s1_write                              : std_logic;                      -- mm_interconnect_0:i2c_sda_s1_write -> mm_interconnect_0_i2c_sda_s1_write:in
	signal mm_interconnect_0_i2c_sda_s1_writedata                          : std_logic_vector(31 downto 0);  -- mm_interconnect_0:i2c_sda_s1_writedata -> i2c_sda:writedata
	signal mm_interconnect_0_sd_cont_0_slave_chipselect                    : std_logic;                      -- mm_interconnect_0:sd_cont_0_slave_chipselect -> sd_cont_0:s_chipselect
	signal mm_interconnect_0_sd_cont_0_slave_readdata                      : std_logic_vector(31 downto 0);  -- sd_cont_0:s_readdata -> mm_interconnect_0:sd_cont_0_slave_readdata
	signal sd_cont_0_slave_waitrequest                                     : std_logic;                      -- sd_cont_0:s_waitrequest_n -> sd_cont_0_slave_waitrequest:in
	signal mm_interconnect_0_sd_cont_0_slave_address                       : std_logic_vector(7 downto 0);   -- mm_interconnect_0:sd_cont_0_slave_address -> sd_cont_0:s_address
	signal mm_interconnect_0_sd_cont_0_slave_read                          : std_logic;                      -- mm_interconnect_0:sd_cont_0_slave_read -> sd_cont_0:s_read
	signal mm_interconnect_0_sd_cont_0_slave_write                         : std_logic;                      -- mm_interconnect_0:sd_cont_0_slave_write -> sd_cont_0:s_write
	signal mm_interconnect_0_sd_cont_0_slave_writedata                     : std_logic_vector(31 downto 0);  -- mm_interconnect_0:sd_cont_0_slave_writedata -> sd_cont_0:s_writedata
	signal mm_interconnect_0_sram_uas_readdata                             : std_logic_vector(15 downto 0);  -- sram:uas_readdata -> mm_interconnect_0:sram_uas_readdata
	signal mm_interconnect_0_sram_uas_waitrequest                          : std_logic;                      -- sram:uas_waitrequest -> mm_interconnect_0:sram_uas_waitrequest
	signal mm_interconnect_0_sram_uas_debugaccess                          : std_logic;                      -- mm_interconnect_0:sram_uas_debugaccess -> sram:uas_debugaccess
	signal mm_interconnect_0_sram_uas_address                              : std_logic_vector(18 downto 0);  -- mm_interconnect_0:sram_uas_address -> sram:uas_address
	signal mm_interconnect_0_sram_uas_read                                 : std_logic;                      -- mm_interconnect_0:sram_uas_read -> sram:uas_read
	signal mm_interconnect_0_sram_uas_byteenable                           : std_logic_vector(1 downto 0);   -- mm_interconnect_0:sram_uas_byteenable -> sram:uas_byteenable
	signal mm_interconnect_0_sram_uas_readdatavalid                        : std_logic;                      -- sram:uas_readdatavalid -> mm_interconnect_0:sram_uas_readdatavalid
	signal mm_interconnect_0_sram_uas_lock                                 : std_logic;                      -- mm_interconnect_0:sram_uas_lock -> sram:uas_lock
	signal mm_interconnect_0_sram_uas_write                                : std_logic;                      -- mm_interconnect_0:sram_uas_write -> sram:uas_write
	signal mm_interconnect_0_sram_uas_writedata                            : std_logic_vector(15 downto 0);  -- mm_interconnect_0:sram_uas_writedata -> sram:uas_writedata
	signal mm_interconnect_0_sram_uas_burstcount                           : std_logic_vector(1 downto 0);   -- mm_interconnect_0:sram_uas_burstcount -> sram:uas_burstcount
	signal mm_interconnect_0_cpu_2_debug_mem_slave_readdata                : std_logic_vector(31 downto 0);  -- cpu_2:debug_mem_slave_readdata -> mm_interconnect_0:cpu_2_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_2_debug_mem_slave_waitrequest             : std_logic;                      -- cpu_2:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_2_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_2_debug_mem_slave_debugaccess             : std_logic;                      -- mm_interconnect_0:cpu_2_debug_mem_slave_debugaccess -> cpu_2:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_2_debug_mem_slave_address                 : std_logic_vector(8 downto 0);   -- mm_interconnect_0:cpu_2_debug_mem_slave_address -> cpu_2:debug_mem_slave_address
	signal mm_interconnect_0_cpu_2_debug_mem_slave_read                    : std_logic;                      -- mm_interconnect_0:cpu_2_debug_mem_slave_read -> cpu_2:debug_mem_slave_read
	signal mm_interconnect_0_cpu_2_debug_mem_slave_byteenable              : std_logic_vector(3 downto 0);   -- mm_interconnect_0:cpu_2_debug_mem_slave_byteenable -> cpu_2:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_2_debug_mem_slave_write                   : std_logic;                      -- mm_interconnect_0:cpu_2_debug_mem_slave_write -> cpu_2:debug_mem_slave_write
	signal mm_interconnect_0_cpu_2_debug_mem_slave_writedata               : std_logic_vector(31 downto 0);  -- mm_interconnect_0:cpu_2_debug_mem_slave_writedata -> cpu_2:debug_mem_slave_writedata
	signal mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_chipselect      : std_logic;                      -- mm_interconnect_0:jtag_uart_2_avalon_jtag_slave_chipselect -> jtag_uart_2:av_chipselect
	signal mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0);  -- jtag_uart_2:av_readdata -> mm_interconnect_0:jtag_uart_2_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_waitrequest     : std_logic;                      -- jtag_uart_2:av_waitrequest -> mm_interconnect_0:jtag_uart_2_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);   -- mm_interconnect_0:jtag_uart_2_avalon_jtag_slave_address -> jtag_uart_2:av_address
	signal mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_read            : std_logic;                      -- mm_interconnect_0:jtag_uart_2_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_write           : std_logic;                      -- mm_interconnect_0:jtag_uart_2_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0);  -- mm_interconnect_0:jtag_uart_2_avalon_jtag_slave_writedata -> jtag_uart_2:av_writedata
	signal mm_interconnect_0_mailbox_simple_3_avmm_msg_receiver_readdata   : std_logic_vector(31 downto 0);  -- mailbox_simple_3:avmm_rcv_readdata -> mm_interconnect_0:mailbox_simple_3_avmm_msg_receiver_readdata
	signal mm_interconnect_0_mailbox_simple_3_avmm_msg_receiver_address    : std_logic_vector(1 downto 0);   -- mm_interconnect_0:mailbox_simple_3_avmm_msg_receiver_address -> mailbox_simple_3:avmm_rcv_address
	signal mm_interconnect_0_mailbox_simple_3_avmm_msg_receiver_read       : std_logic;                      -- mm_interconnect_0:mailbox_simple_3_avmm_msg_receiver_read -> mailbox_simple_3:avmm_rcv_read
	signal mm_interconnect_0_mailbox_simple_3_avmm_msg_receiver_write      : std_logic;                      -- mm_interconnect_0:mailbox_simple_3_avmm_msg_receiver_write -> mailbox_simple_3:avmm_rcv_write
	signal mm_interconnect_0_mailbox_simple_3_avmm_msg_receiver_writedata  : std_logic_vector(31 downto 0);  -- mm_interconnect_0:mailbox_simple_3_avmm_msg_receiver_writedata -> mailbox_simple_3:avmm_rcv_writedata
	signal mm_interconnect_0_mailbox_simple_2_avmm_msg_sender_readdata     : std_logic_vector(31 downto 0);  -- mailbox_simple_2:avmm_snd_readdata -> mm_interconnect_0:mailbox_simple_2_avmm_msg_sender_readdata
	signal mm_interconnect_0_mailbox_simple_2_avmm_msg_sender_waitrequest  : std_logic;                      -- mailbox_simple_2:avmm_snd_waitrequest -> mm_interconnect_0:mailbox_simple_2_avmm_msg_sender_waitrequest
	signal mm_interconnect_0_mailbox_simple_2_avmm_msg_sender_address      : std_logic_vector(1 downto 0);   -- mm_interconnect_0:mailbox_simple_2_avmm_msg_sender_address -> mailbox_simple_2:avmm_snd_address
	signal mm_interconnect_0_mailbox_simple_2_avmm_msg_sender_read         : std_logic;                      -- mm_interconnect_0:mailbox_simple_2_avmm_msg_sender_read -> mailbox_simple_2:avmm_snd_read
	signal mm_interconnect_0_mailbox_simple_2_avmm_msg_sender_write        : std_logic;                      -- mm_interconnect_0:mailbox_simple_2_avmm_msg_sender_write -> mailbox_simple_2:avmm_snd_write
	signal mm_interconnect_0_mailbox_simple_2_avmm_msg_sender_writedata    : std_logic_vector(31 downto 0);  -- mm_interconnect_0:mailbox_simple_2_avmm_msg_sender_writedata -> mailbox_simple_2:avmm_snd_writedata
	signal mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_chipselect      : std_logic;                      -- mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_chipselect -> jtag_uart_1:av_chipselect
	signal mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0);  -- jtag_uart_1:av_readdata -> mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_waitrequest     : std_logic;                      -- jtag_uart_1:av_waitrequest -> mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);   -- mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_address -> jtag_uart_1:av_address
	signal mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read            : std_logic;                      -- mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write           : std_logic;                      -- mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0);  -- mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_writedata -> jtag_uart_1:av_writedata
	signal mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_readdata   : std_logic_vector(31 downto 0);  -- mailbox_simple_0:avmm_rcv_readdata -> mm_interconnect_0:mailbox_simple_0_avmm_msg_receiver_readdata
	signal mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_address    : std_logic_vector(1 downto 0);   -- mm_interconnect_0:mailbox_simple_0_avmm_msg_receiver_address -> mailbox_simple_0:avmm_rcv_address
	signal mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_read       : std_logic;                      -- mm_interconnect_0:mailbox_simple_0_avmm_msg_receiver_read -> mailbox_simple_0:avmm_rcv_read
	signal mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_write      : std_logic;                      -- mm_interconnect_0:mailbox_simple_0_avmm_msg_receiver_write -> mailbox_simple_0:avmm_rcv_write
	signal mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_writedata  : std_logic_vector(31 downto 0);  -- mm_interconnect_0:mailbox_simple_0_avmm_msg_receiver_writedata -> mailbox_simple_0:avmm_rcv_writedata
	signal mm_interconnect_0_mailbox_simple_1_avmm_msg_sender_readdata     : std_logic_vector(31 downto 0);  -- mailbox_simple_1:avmm_snd_readdata -> mm_interconnect_0:mailbox_simple_1_avmm_msg_sender_readdata
	signal mm_interconnect_0_mailbox_simple_1_avmm_msg_sender_waitrequest  : std_logic;                      -- mailbox_simple_1:avmm_snd_waitrequest -> mm_interconnect_0:mailbox_simple_1_avmm_msg_sender_waitrequest
	signal mm_interconnect_0_mailbox_simple_1_avmm_msg_sender_address      : std_logic_vector(1 downto 0);   -- mm_interconnect_0:mailbox_simple_1_avmm_msg_sender_address -> mailbox_simple_1:avmm_snd_address
	signal mm_interconnect_0_mailbox_simple_1_avmm_msg_sender_read         : std_logic;                      -- mm_interconnect_0:mailbox_simple_1_avmm_msg_sender_read -> mailbox_simple_1:avmm_snd_read
	signal mm_interconnect_0_mailbox_simple_1_avmm_msg_sender_write        : std_logic;                      -- mm_interconnect_0:mailbox_simple_1_avmm_msg_sender_write -> mailbox_simple_1:avmm_snd_write
	signal mm_interconnect_0_mailbox_simple_1_avmm_msg_sender_writedata    : std_logic_vector(31 downto 0);  -- mm_interconnect_0:mailbox_simple_1_avmm_msg_sender_writedata -> mailbox_simple_1:avmm_snd_writedata
	signal mm_interconnect_0_cpu_1_debug_mem_slave_readdata                : std_logic_vector(31 downto 0);  -- cpu_1:debug_mem_slave_readdata -> mm_interconnect_0:cpu_1_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_1_debug_mem_slave_waitrequest             : std_logic;                      -- cpu_1:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_1_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_1_debug_mem_slave_debugaccess             : std_logic;                      -- mm_interconnect_0:cpu_1_debug_mem_slave_debugaccess -> cpu_1:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_1_debug_mem_slave_address                 : std_logic_vector(8 downto 0);   -- mm_interconnect_0:cpu_1_debug_mem_slave_address -> cpu_1:debug_mem_slave_address
	signal mm_interconnect_0_cpu_1_debug_mem_slave_read                    : std_logic;                      -- mm_interconnect_0:cpu_1_debug_mem_slave_read -> cpu_1:debug_mem_slave_read
	signal mm_interconnect_0_cpu_1_debug_mem_slave_byteenable              : std_logic_vector(3 downto 0);   -- mm_interconnect_0:cpu_1_debug_mem_slave_byteenable -> cpu_1:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_1_debug_mem_slave_write                   : std_logic;                      -- mm_interconnect_0:cpu_1_debug_mem_slave_write -> cpu_1:debug_mem_slave_write
	signal mm_interconnect_0_cpu_1_debug_mem_slave_writedata               : std_logic_vector(31 downto 0);  -- mm_interconnect_0:cpu_1_debug_mem_slave_writedata -> cpu_1:debug_mem_slave_writedata
	signal video_dma_mm_read_readdata                                      : std_logic_vector(31 downto 0);  -- mm_interconnect_1:video_dma_mm_read_readdata -> video_dma:mm_read_readdata
	signal video_dma_mm_read_waitrequest                                   : std_logic;                      -- mm_interconnect_1:video_dma_mm_read_waitrequest -> video_dma:mm_read_waitrequest
	signal video_dma_mm_read_address                                       : std_logic_vector(28 downto 0);  -- video_dma:mm_read_address -> mm_interconnect_1:video_dma_mm_read_address
	signal video_dma_mm_read_read                                          : std_logic;                      -- video_dma:mm_read_read -> mm_interconnect_1:video_dma_mm_read_read
	signal video_dma_mm_read_byteenable                                    : std_logic_vector(3 downto 0);   -- video_dma:mm_read_byteenable -> mm_interconnect_1:video_dma_mm_read_byteenable
	signal video_dma_mm_read_readdatavalid                                 : std_logic;                      -- mm_interconnect_1:video_dma_mm_read_readdatavalid -> video_dma:mm_read_readdatavalid
	signal video_dma_mm_read_burstcount                                    : std_logic_vector(7 downto 0);   -- video_dma:mm_read_burstcount -> mm_interconnect_1:video_dma_mm_read_burstcount
	signal read_dma_0_mm_read_readdata                                     : std_logic_vector(31 downto 0);  -- mm_interconnect_1:read_dma_0_mm_read_readdata -> read_dma_0:mm_read_readdata
	signal read_dma_0_mm_read_waitrequest                                  : std_logic;                      -- mm_interconnect_1:read_dma_0_mm_read_waitrequest -> read_dma_0:mm_read_waitrequest
	signal read_dma_0_mm_read_address                                      : std_logic_vector(28 downto 0);  -- read_dma_0:mm_read_address -> mm_interconnect_1:read_dma_0_mm_read_address
	signal read_dma_0_mm_read_read                                         : std_logic;                      -- read_dma_0:mm_read_read -> mm_interconnect_1:read_dma_0_mm_read_read
	signal read_dma_0_mm_read_byteenable                                   : std_logic_vector(3 downto 0);   -- read_dma_0:mm_read_byteenable -> mm_interconnect_1:read_dma_0_mm_read_byteenable
	signal read_dma_0_mm_read_readdatavalid                                : std_logic;                      -- mm_interconnect_1:read_dma_0_mm_read_readdatavalid -> read_dma_0:mm_read_readdatavalid
	signal read_dma_0_mm_read_burstcount                                   : std_logic_vector(7 downto 0);   -- read_dma_0:mm_read_burstcount -> mm_interconnect_1:read_dma_0_mm_read_burstcount
	signal mm_interconnect_1_lpddr2_avl_1_beginbursttransfer               : std_logic;                      -- mm_interconnect_1:lpddr2_avl_1_beginbursttransfer -> lpddr2:avl_burstbegin_1
	signal mm_interconnect_1_lpddr2_avl_1_readdata                         : std_logic_vector(31 downto 0);  -- lpddr2:avl_rdata_1 -> mm_interconnect_1:lpddr2_avl_1_readdata
	signal lpddr2_avl_1_waitrequest                                        : std_logic;                      -- lpddr2:avl_ready_1 -> lpddr2_avl_1_waitrequest:in
	signal mm_interconnect_1_lpddr2_avl_1_address                          : std_logic_vector(26 downto 0);  -- mm_interconnect_1:lpddr2_avl_1_address -> lpddr2:avl_addr_1
	signal mm_interconnect_1_lpddr2_avl_1_read                             : std_logic;                      -- mm_interconnect_1:lpddr2_avl_1_read -> lpddr2:avl_read_req_1
	signal mm_interconnect_1_lpddr2_avl_1_byteenable                       : std_logic_vector(3 downto 0);   -- mm_interconnect_1:lpddr2_avl_1_byteenable -> lpddr2:avl_be_1
	signal mm_interconnect_1_lpddr2_avl_1_readdatavalid                    : std_logic;                      -- lpddr2:avl_rdata_valid_1 -> mm_interconnect_1:lpddr2_avl_1_readdatavalid
	signal mm_interconnect_1_lpddr2_avl_1_write                            : std_logic;                      -- mm_interconnect_1:lpddr2_avl_1_write -> lpddr2:avl_write_req_1
	signal mm_interconnect_1_lpddr2_avl_1_writedata                        : std_logic_vector(31 downto 0);  -- mm_interconnect_1:lpddr2_avl_1_writedata -> lpddr2:avl_wdata_1
	signal mm_interconnect_1_lpddr2_avl_1_burstcount                       : std_logic_vector(7 downto 0);   -- mm_interconnect_1:lpddr2_avl_1_burstcount -> lpddr2:avl_size_1
	signal write_dma_0_mm_write_waitrequest                                : std_logic;                      -- mm_interconnect_2:write_dma_0_mm_write_waitrequest -> write_dma_0:mm_write_waitrequest
	signal write_dma_0_mm_write_address                                    : std_logic_vector(28 downto 0);  -- write_dma_0:mm_write_address -> mm_interconnect_2:write_dma_0_mm_write_address
	signal write_dma_0_mm_write_byteenable                                 : std_logic_vector(3 downto 0);   -- write_dma_0:mm_write_byteenable -> mm_interconnect_2:write_dma_0_mm_write_byteenable
	signal write_dma_0_mm_write_write                                      : std_logic;                      -- write_dma_0:mm_write_write -> mm_interconnect_2:write_dma_0_mm_write_write
	signal write_dma_0_mm_write_writedata                                  : std_logic_vector(31 downto 0);  -- write_dma_0:mm_write_writedata -> mm_interconnect_2:write_dma_0_mm_write_writedata
	signal write_dma_0_mm_write_burstcount                                 : std_logic_vector(7 downto 0);   -- write_dma_0:mm_write_burstcount -> mm_interconnect_2:write_dma_0_mm_write_burstcount
	signal mm_interconnect_2_lpddr2_avl_2_beginbursttransfer               : std_logic;                      -- mm_interconnect_2:lpddr2_avl_2_beginbursttransfer -> lpddr2:avl_burstbegin_2
	signal mm_interconnect_2_lpddr2_avl_2_readdata                         : std_logic_vector(31 downto 0);  -- lpddr2:avl_rdata_2 -> mm_interconnect_2:lpddr2_avl_2_readdata
	signal lpddr2_avl_2_waitrequest                                        : std_logic;                      -- lpddr2:avl_ready_2 -> lpddr2_avl_2_waitrequest:in
	signal mm_interconnect_2_lpddr2_avl_2_address                          : std_logic_vector(26 downto 0);  -- mm_interconnect_2:lpddr2_avl_2_address -> lpddr2:avl_addr_2
	signal mm_interconnect_2_lpddr2_avl_2_read                             : std_logic;                      -- mm_interconnect_2:lpddr2_avl_2_read -> lpddr2:avl_read_req_2
	signal mm_interconnect_2_lpddr2_avl_2_byteenable                       : std_logic_vector(3 downto 0);   -- mm_interconnect_2:lpddr2_avl_2_byteenable -> lpddr2:avl_be_2
	signal mm_interconnect_2_lpddr2_avl_2_readdatavalid                    : std_logic;                      -- lpddr2:avl_rdata_valid_2 -> mm_interconnect_2:lpddr2_avl_2_readdatavalid
	signal mm_interconnect_2_lpddr2_avl_2_write                            : std_logic;                      -- mm_interconnect_2:lpddr2_avl_2_write -> lpddr2:avl_write_req_2
	signal mm_interconnect_2_lpddr2_avl_2_writedata                        : std_logic_vector(31 downto 0);  -- mm_interconnect_2:lpddr2_avl_2_writedata -> lpddr2:avl_wdata_2
	signal mm_interconnect_2_lpddr2_avl_2_burstcount                       : std_logic_vector(7 downto 0);   -- mm_interconnect_2:lpddr2_avl_2_burstcount -> lpddr2:avl_size_2
	signal irq_mapper_receiver0_irq                                        : std_logic;                      -- video_dma:csr_irq_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                        : std_logic;                      -- write_dma_0:csr_irq_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                        : std_logic;                      -- read_dma_0:csr_irq_irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                        : std_logic;                      -- mailbox_simple_1:irq_msg -> irq_mapper:receiver3_irq
	signal irq_mapper_receiver4_irq                                        : std_logic;                      -- mailbox_simple_2:irq_msg -> irq_mapper:receiver4_irq
	signal irq_mapper_receiver5_irq                                        : std_logic;                      -- timer_0:irq -> irq_mapper:receiver5_irq
	signal irq_mapper_receiver6_irq                                        : std_logic;                      -- jtag_uart_0:av_irq -> irq_mapper:receiver6_irq
	signal irq_mapper_receiver7_irq                                        : std_logic;                      -- key:irq -> irq_mapper:receiver7_irq
	signal irq_mapper_receiver8_irq                                        : std_logic;                      -- timer_1:irq -> irq_mapper:receiver8_irq
	signal cpu_0_irq_irq                                                   : std_logic_vector(31 downto 0);  -- irq_mapper:sender_irq -> cpu_0:irq
	signal irq_mapper_001_receiver0_irq                                    : std_logic;                      -- mailbox_simple_0:irq_msg -> irq_mapper_001:receiver0_irq
	signal irq_mapper_001_receiver1_irq                                    : std_logic;                      -- jtag_uart_1:av_irq -> irq_mapper_001:receiver1_irq
	signal cpu_1_irq_irq                                                   : std_logic_vector(31 downto 0);  -- irq_mapper_001:sender_irq -> cpu_1:irq
	signal irq_mapper_002_receiver0_irq                                    : std_logic;                      -- mailbox_simple_3:irq_msg -> irq_mapper_002:receiver0_irq
	signal irq_mapper_002_receiver1_irq                                    : std_logic;                      -- jtag_uart_2:av_irq -> irq_mapper_002:receiver1_irq
	signal cpu_2_irq_irq                                                   : std_logic_vector(31 downto 0);  -- irq_mapper_002:sender_irq -> cpu_2:irq
	signal video_fifo_out_valid                                            : std_logic;                      -- video_fifo:avalonst_source_valid -> avalon_st_adapter:in_0_valid
	signal video_fifo_out_data                                             : std_logic_vector(31 downto 0);  -- video_fifo:avalonst_source_data -> avalon_st_adapter:in_0_data
	signal video_fifo_out_ready                                            : std_logic;                      -- avalon_st_adapter:in_0_ready -> video_fifo:avalonst_source_ready
	signal video_fifo_out_startofpacket                                    : std_logic;                      -- video_fifo:avalonst_source_startofpacket -> avalon_st_adapter:in_0_startofpacket
	signal video_fifo_out_endofpacket                                      : std_logic;                      -- video_fifo:avalonst_source_endofpacket -> avalon_st_adapter:in_0_endofpacket
	signal video_fifo_out_empty                                            : std_logic_vector(1 downto 0);   -- video_fifo:avalonst_source_empty -> avalon_st_adapter:in_0_empty
	signal avalon_st_adapter_out_0_valid                                   : std_logic;                      -- avalon_st_adapter:out_0_valid -> Pixel_Con:valid_in
	signal avalon_st_adapter_out_0_data                                    : std_logic_vector(31 downto 0);  -- avalon_st_adapter:out_0_data -> Pixel_Con:data_in
	signal avalon_st_adapter_out_0_ready                                   : std_logic;                      -- Pixel_Con:ready_out -> avalon_st_adapter:out_0_ready
	signal avalon_st_adapter_out_0_startofpacket                           : std_logic;                      -- avalon_st_adapter:out_0_startofpacket -> Pixel_Con:sop_in
	signal avalon_st_adapter_out_0_endofpacket                             : std_logic;                      -- avalon_st_adapter:out_0_endofpacket -> Pixel_Con:eop_in
	signal avalon_st_adapter_out_0_empty                                   : std_logic_vector(1 downto 0);   -- avalon_st_adapter:out_0_empty -> Pixel_Con:empty_in
	signal video_dma_st_source_valid                                       : std_logic;                      -- video_dma:st_source_valid -> avalon_st_adapter_001:in_0_valid
	signal video_dma_st_source_data                                        : std_logic_vector(31 downto 0);  -- video_dma:st_source_data -> avalon_st_adapter_001:in_0_data
	signal video_dma_st_source_ready                                       : std_logic;                      -- avalon_st_adapter_001:in_0_ready -> video_dma:st_source_ready
	signal video_dma_st_source_startofpacket                               : std_logic;                      -- video_dma:st_source_startofpacket -> avalon_st_adapter_001:in_0_startofpacket
	signal video_dma_st_source_endofpacket                                 : std_logic;                      -- video_dma:st_source_endofpacket -> avalon_st_adapter_001:in_0_endofpacket
	signal video_dma_st_source_empty                                       : std_logic_vector(1 downto 0);   -- video_dma:st_source_empty -> avalon_st_adapter_001:in_0_empty
	signal avalon_st_adapter_001_out_0_valid                               : std_logic;                      -- avalon_st_adapter_001:out_0_valid -> video_fifo:avalonst_sink_valid
	signal avalon_st_adapter_001_out_0_data                                : std_logic_vector(31 downto 0);  -- avalon_st_adapter_001:out_0_data -> video_fifo:avalonst_sink_data
	signal avalon_st_adapter_001_out_0_ready                               : std_logic;                      -- video_fifo:avalonst_sink_ready -> avalon_st_adapter_001:out_0_ready
	signal avalon_st_adapter_001_out_0_startofpacket                       : std_logic;                      -- avalon_st_adapter_001:out_0_startofpacket -> video_fifo:avalonst_sink_startofpacket
	signal avalon_st_adapter_001_out_0_endofpacket                         : std_logic;                      -- avalon_st_adapter_001:out_0_endofpacket -> video_fifo:avalonst_sink_endofpacket
	signal avalon_st_adapter_001_out_0_empty                               : std_logic_vector(1 downto 0);   -- avalon_st_adapter_001:out_0_empty -> video_fifo:avalonst_sink_empty
	signal rst_controller_reset_out_reset                                  : std_logic;                      -- rst_controller:reset_out -> [avalon_st_adapter:in_rst_0_reset, rst_controller_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset                              : std_logic;                      -- rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:cpu_0_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_001_reset_out_reset_req                          : std_logic;                      -- rst_controller_001:reset_req -> [cpu_0:reset_req, rst_translator:reset_req_in]
	signal cpu_0_debug_reset_request_reset                                 : std_logic;                      -- cpu_0:debug_reset_request -> rst_controller_001:reset_in0
	signal rst_controller_002_reset_out_reset                              : std_logic;                      -- rst_controller_002:reset_out -> [irq_mapper_001:reset, mm_interconnect_0:cpu_1_reset_reset_bridge_in_reset_reset, rst_controller_002_reset_out_reset:in, rst_translator_001:in_reset]
	signal rst_controller_002_reset_out_reset_req                          : std_logic;                      -- rst_controller_002:reset_req -> [cpu_1:reset_req, rst_translator_001:reset_req_in]
	signal cpu_1_debug_reset_request_reset                                 : std_logic;                      -- cpu_1:debug_reset_request -> rst_controller_002:reset_in0
	signal rst_controller_003_reset_out_reset                              : std_logic;                      -- rst_controller_003:reset_out -> [irq_mapper_002:reset, mm_interconnect_0:cpu_2_reset_reset_bridge_in_reset_reset, rst_controller_003_reset_out_reset:in, rst_translator_002:in_reset]
	signal rst_controller_003_reset_out_reset_req                          : std_logic;                      -- rst_controller_003:reset_req -> [cpu_2:reset_req, rst_translator_002:reset_req_in]
	signal cpu_2_debug_reset_request_reset                                 : std_logic;                      -- cpu_2:debug_reset_request -> rst_controller_003:reset_in0
	signal rst_controller_004_reset_out_reset                              : std_logic;                      -- rst_controller_004:reset_out -> [avalon_st_adapter_001:in_rst_0_reset, mm_interconnect_0:lpddr2_mp_cmd_reset_n_0_reset_bridge_in_reset_reset, mm_interconnect_0:mailbox_simple_1_rst_n_reset_bridge_in_reset_reset, mm_interconnect_1:lpddr2_mp_cmd_reset_n_1_reset_bridge_in_reset_reset, mm_interconnect_1:video_dma_reset_n_reset_bridge_in_reset_reset, mm_interconnect_2:lpddr2_mp_cmd_reset_n_2_reset_bridge_in_reset_reset, mm_interconnect_2:write_dma_0_reset_n_reset_bridge_in_reset_reset, rst_controller_004_reset_out_reset:in, sram:reset_reset, sram_bridge:reset, sram_sharer:reset_reset, twod_idct_st_hw_0:reset]
	signal rst_controller_005_reset_out_reset                              : std_logic;                      -- rst_controller_005:reset_out -> [mm_interconnect_0:sd_cont_0_reset_reset_bridge_in_reset_reset, sd_cont_0:reset]
	signal reset_reset_n_ports_inv                                         : std_logic;                      -- reset_reset_n:inv -> reset_controller_0:reset_in0
	signal reset_controller_0_reset_out_reset_ports_inv                    : std_logic;                      -- reset_controller_0_reset_out_reset:inv -> [lpddr2:mp_cmd_reset_n_0_reset_n, lpddr2:mp_cmd_reset_n_1_reset_n, lpddr2:mp_cmd_reset_n_2_reset_n, lpddr2:mp_rfifo_reset_n_0_reset_n, lpddr2:mp_rfifo_reset_n_1_reset_n, lpddr2:mp_wfifo_reset_n_0_reset_n, lpddr2:mp_wfifo_reset_n_1_reset_n, lpddr2:soft_reset_n]
	signal sd_cont_0_master_inv                                            : std_logic;                      -- mm_interconnect_0_sd_cont_0_master_waitrequest:inv -> sd_cont_0:m_waitrequest_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv  : std_logic;                      -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv : std_logic;                      -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_lpddr2_avl_0_inv                              : std_logic;                      -- lpddr2_avl_0_waitrequest:inv -> mm_interconnect_0:lpddr2_avl_0_waitrequest
	signal mm_interconnect_0_timer_0_s1_write_ports_inv                    : std_logic;                      -- mm_interconnect_0_timer_0_s1_write:inv -> timer_0:write_n
	signal mm_interconnect_0_key_s1_write_ports_inv                        : std_logic;                      -- mm_interconnect_0_key_s1_write:inv -> key:write_n
	signal mm_interconnect_0_timer_1_s1_write_ports_inv                    : std_logic;                      -- mm_interconnect_0_timer_1_s1_write:inv -> timer_1:write_n
	signal mm_interconnect_0_ledg_s1_write_ports_inv                       : std_logic;                      -- mm_interconnect_0_ledg_s1_write:inv -> ledg:write_n
	signal mm_interconnect_0_ledr_s1_write_ports_inv                       : std_logic;                      -- mm_interconnect_0_ledr_s1_write:inv -> ledr:write_n
	signal mm_interconnect_0_i2c_scl_s1_write_ports_inv                    : std_logic;                      -- mm_interconnect_0_i2c_scl_s1_write:inv -> i2c_scl:write_n
	signal mm_interconnect_0_i2c_sda_s1_write_ports_inv                    : std_logic;                      -- mm_interconnect_0_i2c_sda_s1_write:inv -> i2c_sda:write_n
	signal mm_interconnect_0_sd_cont_0_slave_inv                           : std_logic;                      -- sd_cont_0_slave_waitrequest:inv -> mm_interconnect_0:sd_cont_0_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_read_ports_inv  : std_logic;                      -- mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_read:inv -> jtag_uart_2:av_read_n
	signal mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_write_ports_inv : std_logic;                      -- mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_write:inv -> jtag_uart_2:av_write_n
	signal mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read_ports_inv  : std_logic;                      -- mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read:inv -> jtag_uart_1:av_read_n
	signal mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write_ports_inv : std_logic;                      -- mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write:inv -> jtag_uart_1:av_write_n
	signal mm_interconnect_1_lpddr2_avl_1_inv                              : std_logic;                      -- lpddr2_avl_1_waitrequest:inv -> mm_interconnect_1:lpddr2_avl_1_waitrequest
	signal mm_interconnect_2_lpddr2_avl_2_inv                              : std_logic;                      -- lpddr2_avl_2_waitrequest:inv -> mm_interconnect_2:lpddr2_avl_2_waitrequest
	signal rst_controller_reset_out_reset_ports_inv                        : std_logic;                      -- rst_controller_reset_out_reset:inv -> [Pixel_Con:reset_n, video:reset_n, video_fifo:rdreset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                    : std_logic;                      -- rst_controller_001_reset_out_reset:inv -> [cpu_0:reset_n, jtag_uart_0:rst_n]
	signal rst_controller_002_reset_out_reset_ports_inv                    : std_logic;                      -- rst_controller_002_reset_out_reset:inv -> [cpu_1:reset_n, jtag_uart_1:rst_n]
	signal rst_controller_003_reset_out_reset_ports_inv                    : std_logic;                      -- rst_controller_003_reset_out_reset:inv -> [cpu_2:reset_n, jtag_uart_2:rst_n]
	signal rst_controller_004_reset_out_reset_ports_inv                    : std_logic;                      -- rst_controller_004_reset_out_reset:inv -> [i2c_scl:reset_n, i2c_sda:reset_n, key:reset_n, ledg:reset_n, ledr:reset_n, mailbox_simple_0:rst_n, mailbox_simple_1:rst_n, mailbox_simple_2:rst_n, mailbox_simple_3:rst_n, read_dma_0:reset_n_reset_n, sysid:reset_n, timer_0:reset_n, timer_1:reset_n, video_dma:reset_n_reset_n, video_fifo:wrreset_n, write_dma_0:reset_n_reset_n]

begin

	pixel_con : component Pixel_Conv
		generic map (
			SOURCE_SYMBOLS_PER_BEAT => 1
		)
		port map (
			clk       => video_pll_outclk0_clk,                    --       clk.clk
			reset_n   => rst_controller_reset_out_reset_ports_inv, -- clk_reset.reset_n
			ready_out => avalon_st_adapter_out_0_ready,            --        in.ready
			valid_in  => avalon_st_adapter_out_0_valid,            --          .valid
			data_in   => avalon_st_adapter_out_0_data,             --          .data
			eop_in    => avalon_st_adapter_out_0_endofpacket,      --          .endofpacket
			sop_in    => avalon_st_adapter_out_0_startofpacket,    --          .startofpacket
			empty_in  => avalon_st_adapter_out_0_empty,            --          .empty
			ready_in  => pixel_con_out_ready,                      --       out.ready
			valid_out => pixel_con_out_valid,                      --          .valid
			data_out  => pixel_con_out_data,                       --          .data
			eop_out   => pixel_con_out_endofpacket,                --          .endofpacket
			sop_out   => pixel_con_out_startofpacket,              --          .startofpacket
			empty_out => pixel_con_out_empty                       --          .empty
		);

	cpu_0 : component HW_QSYS_cpu_0
		port map (
			clk                                 => clk_125_clk,                                         --                       clk.clk
			reset_n                             => rst_controller_001_reset_out_reset_ports_inv,        --                     reset.reset_n
			reset_req                           => rst_controller_001_reset_out_reset_req,              --                          .reset_req
			d_address                           => cpu_0_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_0_data_master_read,                              --                          .read
			d_readdata                          => cpu_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_0_data_master_write,                             --                          .write
			d_writedata                         => cpu_0_data_master_writedata,                         --                          .writedata
			d_burstcount                        => cpu_0_data_master_burstcount,                        --                          .burstcount
			d_readdatavalid                     => cpu_0_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => cpu_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_0_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_0_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => cpu_0_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => cpu_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                 -- custom_instruction_master.readra
		);

	cpu_1 : component HW_QSYS_cpu_1
		port map (
			clk                                 => clk_125_clk,                                         --                       clk.clk
			reset_n                             => rst_controller_002_reset_out_reset_ports_inv,        --                     reset.reset_n
			reset_req                           => rst_controller_002_reset_out_reset_req,              --                          .reset_req
			d_address                           => cpu_1_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_1_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_1_data_master_read,                              --                          .read
			d_readdata                          => cpu_1_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_1_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_1_data_master_write,                             --                          .write
			d_writedata                         => cpu_1_data_master_writedata,                         --                          .writedata
			d_burstcount                        => cpu_1_data_master_burstcount,                        --                          .burstcount
			d_readdatavalid                     => cpu_1_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => cpu_1_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_1_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_1_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_1_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_1_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => cpu_1_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => cpu_1_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_1_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_1_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_1_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_1_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_1_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_1_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_1_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_1_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_1_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                 -- custom_instruction_master.readra
		);

	cpu_2 : component HW_QSYS_cpu_2
		port map (
			clk                                 => clk_125_clk,                                         --                       clk.clk
			reset_n                             => rst_controller_003_reset_out_reset_ports_inv,        --                     reset.reset_n
			reset_req                           => rst_controller_003_reset_out_reset_req,              --                          .reset_req
			d_address                           => cpu_2_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_2_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_2_data_master_read,                              --                          .read
			d_readdata                          => cpu_2_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_2_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_2_data_master_write,                             --                          .write
			d_writedata                         => cpu_2_data_master_writedata,                         --                          .writedata
			d_burstcount                        => cpu_2_data_master_burstcount,                        --                          .burstcount
			d_readdatavalid                     => cpu_2_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => cpu_2_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_2_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_2_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_2_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_2_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => cpu_2_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => cpu_2_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_2_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_2_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_2_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_2_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_2_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_2_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_2_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_2_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_2_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                 -- custom_instruction_master.readra
		);

	i2c_scl : component HW_QSYS_i2c_scl
		port map (
			clk        => clk_125_clk,                                  --                 clk.clk
			reset_n    => rst_controller_004_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_i2c_scl_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_i2c_scl_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_i2c_scl_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_i2c_scl_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_i2c_scl_s1_readdata,        --                    .readdata
			out_port   => i2c_scl_export                                -- external_connection.export
		);

	i2c_sda : component HW_QSYS_i2c_sda
		port map (
			clk        => clk_125_clk,                                  --                 clk.clk
			reset_n    => rst_controller_004_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_i2c_sda_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_i2c_sda_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_i2c_sda_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_i2c_sda_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_i2c_sda_s1_readdata,        --                    .readdata
			bidir_port => i2c_sda_export                                -- external_connection.export
		);

	jtag_uart_0 : component HW_QSYS_jtag_uart_0
		port map (
			clk            => clk_125_clk,                                                     --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv,                    --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver6_irq                                         --               irq.irq
		);

	jtag_uart_1 : component HW_QSYS_jtag_uart_0
		port map (
			clk            => clk_125_clk,                                                     --               clk.clk
			rst_n          => rst_controller_002_reset_out_reset_ports_inv,                    --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_001_receiver1_irq                                     --               irq.irq
		);

	jtag_uart_2 : component HW_QSYS_jtag_uart_0
		port map (
			clk            => clk_125_clk,                                                     --               clk.clk
			rst_n          => rst_controller_003_reset_out_reset_ports_inv,                    --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_002_receiver1_irq                                     --               irq.irq
		);

	key : component HW_QSYS_key
		port map (
			clk        => clk_125_clk,                                  --                 clk.clk
			reset_n    => rst_controller_004_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_key_s1_address,             --                  s1.address
			write_n    => mm_interconnect_0_key_s1_write_ports_inv,     --                    .write_n
			writedata  => mm_interconnect_0_key_s1_writedata,           --                    .writedata
			chipselect => mm_interconnect_0_key_s1_chipselect,          --                    .chipselect
			readdata   => mm_interconnect_0_key_s1_readdata,            --                    .readdata
			in_port    => key_export,                                   -- external_connection.export
			irq        => irq_mapper_receiver7_irq                      --                 irq.irq
		);

	ledg : component HW_QSYS_ledg
		port map (
			clk        => clk_125_clk,                                  --                 clk.clk
			reset_n    => rst_controller_004_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_ledg_s1_address,            --                  s1.address
			write_n    => mm_interconnect_0_ledg_s1_write_ports_inv,    --                    .write_n
			writedata  => mm_interconnect_0_ledg_s1_writedata,          --                    .writedata
			chipselect => mm_interconnect_0_ledg_s1_chipselect,         --                    .chipselect
			readdata   => mm_interconnect_0_ledg_s1_readdata,           --                    .readdata
			out_port   => ledg_export                                   -- external_connection.export
		);

	ledr : component HW_QSYS_ledg
		port map (
			clk        => clk_125_clk,                                  --                 clk.clk
			reset_n    => rst_controller_004_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_ledr_s1_address,            --                  s1.address
			write_n    => mm_interconnect_0_ledr_s1_write_ports_inv,    --                    .write_n
			writedata  => mm_interconnect_0_ledr_s1_writedata,          --                    .writedata
			chipselect => mm_interconnect_0_ledr_s1_chipselect,         --                    .chipselect
			readdata   => mm_interconnect_0_ledr_s1_readdata,           --                    .readdata
			out_port   => ledr_export                                   -- external_connection.export
		);

	lpddr2 : component HW_QSYS_lpddr2
		port map (
			pll_ref_clk                => lpddr2_pll_ref_clk_clk,                            --        pll_ref_clk.clk
			global_reset_n             => lpddr2_global_reset_reset_n,                       --       global_reset.reset_n
			soft_reset_n               => reset_controller_0_reset_out_reset_ports_inv,      --         soft_reset.reset_n
			afi_clk                    => open,                                              --            afi_clk.clk
			afi_half_clk               => open,                                              --       afi_half_clk.clk
			afi_reset_n                => open,                                              --          afi_reset.reset_n
			afi_reset_export_n         => open,                                              --   afi_reset_export.reset_n
			mem_ca                     => lpddr2_mem_ca,                                     --             memory.mem_ca
			mem_ck                     => lpddr2_mem_ck,                                     --                   .mem_ck
			mem_ck_n                   => lpddr2_mem_ck_n,                                   --                   .mem_ck_n
			mem_cke                    => lpddr2_mem_cke,                                    --                   .mem_cke
			mem_cs_n                   => lpddr2_mem_cs_n,                                   --                   .mem_cs_n
			mem_dm                     => lpddr2_mem_dm,                                     --                   .mem_dm
			mem_dq                     => lpddr2_mem_dq,                                     --                   .mem_dq
			mem_dqs                    => lpddr2_mem_dqs,                                    --                   .mem_dqs
			mem_dqs_n                  => lpddr2_mem_dqs_n,                                  --                   .mem_dqs_n
			avl_ready_0                => lpddr2_avl_0_waitrequest,                          --              avl_0.waitrequest_n
			avl_burstbegin_0           => mm_interconnect_0_lpddr2_avl_0_beginbursttransfer, --                   .beginbursttransfer
			avl_addr_0                 => mm_interconnect_0_lpddr2_avl_0_address,            --                   .address
			avl_rdata_valid_0          => mm_interconnect_0_lpddr2_avl_0_readdatavalid,      --                   .readdatavalid
			avl_rdata_0                => mm_interconnect_0_lpddr2_avl_0_readdata,           --                   .readdata
			avl_wdata_0                => mm_interconnect_0_lpddr2_avl_0_writedata,          --                   .writedata
			avl_be_0                   => mm_interconnect_0_lpddr2_avl_0_byteenable,         --                   .byteenable
			avl_read_req_0             => mm_interconnect_0_lpddr2_avl_0_read,               --                   .read
			avl_write_req_0            => mm_interconnect_0_lpddr2_avl_0_write,              --                   .write
			avl_size_0                 => mm_interconnect_0_lpddr2_avl_0_burstcount,         --                   .burstcount
			avl_ready_1                => lpddr2_avl_1_waitrequest,                          --              avl_1.waitrequest_n
			avl_burstbegin_1           => mm_interconnect_1_lpddr2_avl_1_beginbursttransfer, --                   .beginbursttransfer
			avl_addr_1                 => mm_interconnect_1_lpddr2_avl_1_address,            --                   .address
			avl_rdata_valid_1          => mm_interconnect_1_lpddr2_avl_1_readdatavalid,      --                   .readdatavalid
			avl_rdata_1                => mm_interconnect_1_lpddr2_avl_1_readdata,           --                   .readdata
			avl_wdata_1                => mm_interconnect_1_lpddr2_avl_1_writedata,          --                   .writedata
			avl_be_1                   => mm_interconnect_1_lpddr2_avl_1_byteenable,         --                   .byteenable
			avl_read_req_1             => mm_interconnect_1_lpddr2_avl_1_read,               --                   .read
			avl_write_req_1            => mm_interconnect_1_lpddr2_avl_1_write,              --                   .write
			avl_size_1                 => mm_interconnect_1_lpddr2_avl_1_burstcount,         --                   .burstcount
			avl_ready_2                => lpddr2_avl_2_waitrequest,                          --              avl_2.waitrequest_n
			avl_burstbegin_2           => mm_interconnect_2_lpddr2_avl_2_beginbursttransfer, --                   .beginbursttransfer
			avl_addr_2                 => mm_interconnect_2_lpddr2_avl_2_address,            --                   .address
			avl_rdata_valid_2          => mm_interconnect_2_lpddr2_avl_2_readdatavalid,      --                   .readdatavalid
			avl_rdata_2                => mm_interconnect_2_lpddr2_avl_2_readdata,           --                   .readdata
			avl_wdata_2                => mm_interconnect_2_lpddr2_avl_2_writedata,          --                   .writedata
			avl_be_2                   => mm_interconnect_2_lpddr2_avl_2_byteenable,         --                   .byteenable
			avl_read_req_2             => mm_interconnect_2_lpddr2_avl_2_read,               --                   .read
			avl_write_req_2            => mm_interconnect_2_lpddr2_avl_2_write,              --                   .write
			avl_size_2                 => mm_interconnect_2_lpddr2_avl_2_burstcount,         --                   .burstcount
			mp_cmd_clk_0_clk           => clk_125_clk,                                       --       mp_cmd_clk_0.clk
			mp_cmd_reset_n_0_reset_n   => reset_controller_0_reset_out_reset_ports_inv,      --   mp_cmd_reset_n_0.reset_n
			mp_cmd_clk_1_clk           => clk_125_clk,                                       --       mp_cmd_clk_1.clk
			mp_cmd_reset_n_1_reset_n   => reset_controller_0_reset_out_reset_ports_inv,      --   mp_cmd_reset_n_1.reset_n
			mp_cmd_clk_2_clk           => clk_125_clk,                                       --       mp_cmd_clk_2.clk
			mp_cmd_reset_n_2_reset_n   => reset_controller_0_reset_out_reset_ports_inv,      --   mp_cmd_reset_n_2.reset_n
			mp_rfifo_clk_0_clk         => clk_125_clk,                                       --     mp_rfifo_clk_0.clk
			mp_rfifo_reset_n_0_reset_n => reset_controller_0_reset_out_reset_ports_inv,      -- mp_rfifo_reset_n_0.reset_n
			mp_wfifo_clk_0_clk         => clk_125_clk,                                       --     mp_wfifo_clk_0.clk
			mp_wfifo_reset_n_0_reset_n => reset_controller_0_reset_out_reset_ports_inv,      -- mp_wfifo_reset_n_0.reset_n
			mp_rfifo_clk_1_clk         => clk_125_clk,                                       --     mp_rfifo_clk_1.clk
			mp_rfifo_reset_n_1_reset_n => reset_controller_0_reset_out_reset_ports_inv,      -- mp_rfifo_reset_n_1.reset_n
			mp_wfifo_clk_1_clk         => clk_125_clk,                                       --     mp_wfifo_clk_1.clk
			mp_wfifo_reset_n_1_reset_n => reset_controller_0_reset_out_reset_ports_inv,      -- mp_wfifo_reset_n_1.reset_n
			local_init_done            => lpddr2_status_local_init_done,                     --             status.local_init_done
			local_cal_success          => lpddr2_status_local_cal_success,                   --                   .local_cal_success
			local_cal_fail             => lpddr2_status_local_cal_fail,                      --                   .local_cal_fail
			oct_rzqin                  => lpddr2_oct_rzqin,                                  --                oct.rzqin
			pll_mem_clk                => lpddr2_pll_sharing_pll_mem_clk,                    --        pll_sharing.pll_mem_clk
			pll_write_clk              => lpddr2_pll_sharing_pll_write_clk,                  --                   .pll_write_clk
			pll_locked                 => lpddr2_pll_sharing_pll_locked,                     --                   .pll_locked
			pll_write_clk_pre_phy_clk  => lpddr2_pll_sharing_pll_write_clk_pre_phy_clk,      --                   .pll_write_clk_pre_phy_clk
			pll_addr_cmd_clk           => lpddr2_pll_sharing_pll_addr_cmd_clk,               --                   .pll_addr_cmd_clk
			pll_avl_clk                => lpddr2_pll_sharing_pll_avl_clk,                    --                   .pll_avl_clk
			pll_config_clk             => lpddr2_pll_sharing_pll_config_clk,                 --                   .pll_config_clk
			pll_mem_phy_clk            => lpddr2_pll_sharing_pll_mem_phy_clk,                --                   .pll_mem_phy_clk
			afi_phy_clk                => lpddr2_pll_sharing_afi_phy_clk,                    --                   .afi_phy_clk
			pll_avl_phy_clk            => lpddr2_pll_sharing_pll_avl_phy_clk                 --                   .pll_avl_phy_clk
		);

	mailbox_simple_0 : component altera_avalon_mailbox
		generic map (
			DWIDTH => 32,
			AWIDTH => 2
		)
		port map (
			clk                  => clk_125_clk,                                                    --                   clk.clk
			rst_n                => rst_controller_004_reset_out_reset_ports_inv,                   --                 rst_n.reset_n
			avmm_snd_address     => mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_address,     --       avmm_msg_sender.address
			avmm_snd_writedata   => mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_writedata,   --                      .writedata
			avmm_snd_write       => mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_write,       --                      .write
			avmm_snd_read        => mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_read,        --                      .read
			avmm_snd_readdata    => mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_readdata,    --                      .readdata
			avmm_snd_waitrequest => mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_waitrequest, --                      .waitrequest
			irq_msg              => irq_mapper_001_receiver0_irq,                                   -- interrupt_msg_pending.irq
			avmm_rcv_address     => mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_address,   --     avmm_msg_receiver.address
			avmm_rcv_read        => mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_read,      --                      .read
			avmm_rcv_writedata   => mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_writedata, --                      .writedata
			avmm_rcv_write       => mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_write,     --                      .write
			avmm_rcv_readdata    => mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_readdata,  --                      .readdata
			irq_space            => open                                                            --           (terminated)
		);

	mailbox_simple_1 : component altera_avalon_mailbox
		generic map (
			DWIDTH => 32,
			AWIDTH => 2
		)
		port map (
			clk                  => clk_125_clk,                                                    --                   clk.clk
			rst_n                => rst_controller_004_reset_out_reset_ports_inv,                   --                 rst_n.reset_n
			avmm_snd_address     => mm_interconnect_0_mailbox_simple_1_avmm_msg_sender_address,     --       avmm_msg_sender.address
			avmm_snd_writedata   => mm_interconnect_0_mailbox_simple_1_avmm_msg_sender_writedata,   --                      .writedata
			avmm_snd_write       => mm_interconnect_0_mailbox_simple_1_avmm_msg_sender_write,       --                      .write
			avmm_snd_read        => mm_interconnect_0_mailbox_simple_1_avmm_msg_sender_read,        --                      .read
			avmm_snd_readdata    => mm_interconnect_0_mailbox_simple_1_avmm_msg_sender_readdata,    --                      .readdata
			avmm_snd_waitrequest => mm_interconnect_0_mailbox_simple_1_avmm_msg_sender_waitrequest, --                      .waitrequest
			irq_msg              => irq_mapper_receiver3_irq,                                       -- interrupt_msg_pending.irq
			avmm_rcv_address     => mm_interconnect_0_mailbox_simple_1_avmm_msg_receiver_address,   --     avmm_msg_receiver.address
			avmm_rcv_read        => mm_interconnect_0_mailbox_simple_1_avmm_msg_receiver_read,      --                      .read
			avmm_rcv_writedata   => mm_interconnect_0_mailbox_simple_1_avmm_msg_receiver_writedata, --                      .writedata
			avmm_rcv_write       => mm_interconnect_0_mailbox_simple_1_avmm_msg_receiver_write,     --                      .write
			avmm_rcv_readdata    => mm_interconnect_0_mailbox_simple_1_avmm_msg_receiver_readdata,  --                      .readdata
			irq_space            => open                                                            --           (terminated)
		);

	mailbox_simple_2 : component altera_avalon_mailbox
		generic map (
			DWIDTH => 32,
			AWIDTH => 2
		)
		port map (
			clk                  => clk_125_clk,                                                    --                   clk.clk
			rst_n                => rst_controller_004_reset_out_reset_ports_inv,                   --                 rst_n.reset_n
			avmm_snd_address     => mm_interconnect_0_mailbox_simple_2_avmm_msg_sender_address,     --       avmm_msg_sender.address
			avmm_snd_writedata   => mm_interconnect_0_mailbox_simple_2_avmm_msg_sender_writedata,   --                      .writedata
			avmm_snd_write       => mm_interconnect_0_mailbox_simple_2_avmm_msg_sender_write,       --                      .write
			avmm_snd_read        => mm_interconnect_0_mailbox_simple_2_avmm_msg_sender_read,        --                      .read
			avmm_snd_readdata    => mm_interconnect_0_mailbox_simple_2_avmm_msg_sender_readdata,    --                      .readdata
			avmm_snd_waitrequest => mm_interconnect_0_mailbox_simple_2_avmm_msg_sender_waitrequest, --                      .waitrequest
			irq_msg              => irq_mapper_receiver4_irq,                                       -- interrupt_msg_pending.irq
			avmm_rcv_address     => mm_interconnect_0_mailbox_simple_2_avmm_msg_receiver_address,   --     avmm_msg_receiver.address
			avmm_rcv_read        => mm_interconnect_0_mailbox_simple_2_avmm_msg_receiver_read,      --                      .read
			avmm_rcv_writedata   => mm_interconnect_0_mailbox_simple_2_avmm_msg_receiver_writedata, --                      .writedata
			avmm_rcv_write       => mm_interconnect_0_mailbox_simple_2_avmm_msg_receiver_write,     --                      .write
			avmm_rcv_readdata    => mm_interconnect_0_mailbox_simple_2_avmm_msg_receiver_readdata,  --                      .readdata
			irq_space            => open                                                            --           (terminated)
		);

	mailbox_simple_3 : component altera_avalon_mailbox
		generic map (
			DWIDTH => 32,
			AWIDTH => 2
		)
		port map (
			clk                  => clk_125_clk,                                                    --                   clk.clk
			rst_n                => rst_controller_004_reset_out_reset_ports_inv,                   --                 rst_n.reset_n
			avmm_snd_address     => mm_interconnect_0_mailbox_simple_3_avmm_msg_sender_address,     --       avmm_msg_sender.address
			avmm_snd_writedata   => mm_interconnect_0_mailbox_simple_3_avmm_msg_sender_writedata,   --                      .writedata
			avmm_snd_write       => mm_interconnect_0_mailbox_simple_3_avmm_msg_sender_write,       --                      .write
			avmm_snd_read        => mm_interconnect_0_mailbox_simple_3_avmm_msg_sender_read,        --                      .read
			avmm_snd_readdata    => mm_interconnect_0_mailbox_simple_3_avmm_msg_sender_readdata,    --                      .readdata
			avmm_snd_waitrequest => mm_interconnect_0_mailbox_simple_3_avmm_msg_sender_waitrequest, --                      .waitrequest
			irq_msg              => irq_mapper_002_receiver0_irq,                                   -- interrupt_msg_pending.irq
			avmm_rcv_address     => mm_interconnect_0_mailbox_simple_3_avmm_msg_receiver_address,   --     avmm_msg_receiver.address
			avmm_rcv_read        => mm_interconnect_0_mailbox_simple_3_avmm_msg_receiver_read,      --                      .read
			avmm_rcv_writedata   => mm_interconnect_0_mailbox_simple_3_avmm_msg_receiver_writedata, --                      .writedata
			avmm_rcv_write       => mm_interconnect_0_mailbox_simple_3_avmm_msg_receiver_write,     --                      .write
			avmm_rcv_readdata    => mm_interconnect_0_mailbox_simple_3_avmm_msg_receiver_readdata,  --                      .readdata
			irq_space            => open                                                            --           (terminated)
		);

	read_dma_0 : component HW_QSYS_read_dma_0
		port map (
			mm_read_address              => read_dma_0_mm_read_address,                                --          mm_read.address
			mm_read_read                 => read_dma_0_mm_read_read,                                   --                 .read
			mm_read_byteenable           => read_dma_0_mm_read_byteenable,                             --                 .byteenable
			mm_read_readdata             => read_dma_0_mm_read_readdata,                               --                 .readdata
			mm_read_waitrequest          => read_dma_0_mm_read_waitrequest,                            --                 .waitrequest
			mm_read_readdatavalid        => read_dma_0_mm_read_readdatavalid,                          --                 .readdatavalid
			mm_read_burstcount           => read_dma_0_mm_read_burstcount,                             --                 .burstcount
			clock_clk                    => clk_125_clk,                                               --            clock.clk
			reset_n_reset_n              => rst_controller_004_reset_out_reset_ports_inv,              --          reset_n.reset_n
			csr_writedata                => mm_interconnect_0_read_dma_0_csr_writedata,                --              csr.writedata
			csr_write                    => mm_interconnect_0_read_dma_0_csr_write,                    --                 .write
			csr_byteenable               => mm_interconnect_0_read_dma_0_csr_byteenable,               --                 .byteenable
			csr_readdata                 => mm_interconnect_0_read_dma_0_csr_readdata,                 --                 .readdata
			csr_read                     => mm_interconnect_0_read_dma_0_csr_read,                     --                 .read
			csr_address                  => mm_interconnect_0_read_dma_0_csr_address,                  --                 .address
			descriptor_slave_write       => mm_interconnect_0_read_dma_0_descriptor_slave_write,       -- descriptor_slave.write
			descriptor_slave_waitrequest => mm_interconnect_0_read_dma_0_descriptor_slave_waitrequest, --                 .waitrequest
			descriptor_slave_writedata   => mm_interconnect_0_read_dma_0_descriptor_slave_writedata,   --                 .writedata
			descriptor_slave_byteenable  => mm_interconnect_0_read_dma_0_descriptor_slave_byteenable,  --                 .byteenable
			csr_irq_irq                  => irq_mapper_receiver2_irq,                                  --          csr_irq.irq
			st_source_data               => read_dma_0_st_source_data,                                 --        st_source.data
			st_source_valid              => read_dma_0_st_source_valid,                                --                 .valid
			st_source_ready              => read_dma_0_st_source_ready                                 --                 .ready
		);

	reset_controller_0 : component HW_qsys_reset_controller_0
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "both",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_125_clk,                        --       clk.clk
			reset_out      => reset_controller_0_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	sd_cont_0 : component sd_cont
		port map (
			clk             => clk_50_clk,                                   --  clock.clk
			reset           => rst_controller_005_reset_out_reset,           --  reset.reset
			s_address       => mm_interconnect_0_sd_cont_0_slave_address,    --  slave.address
			s_read          => mm_interconnect_0_sd_cont_0_slave_read,       --       .read
			s_readdata      => mm_interconnect_0_sd_cont_0_slave_readdata,   --       .readdata
			s_write         => mm_interconnect_0_sd_cont_0_slave_write,      --       .write
			s_writedata     => mm_interconnect_0_sd_cont_0_slave_writedata,  --       .writedata
			s_chipselect    => mm_interconnect_0_sd_cont_0_slave_chipselect, --       .chipselect
			s_waitrequest_n => sd_cont_0_slave_waitrequest,                  --       .waitrequest_n
			m_address       => sd_cont_0_master_address,                     -- master.address
			m_read          => sd_cont_0_master_read,                        --       .read
			m_readdata      => sd_cont_0_master_readdata,                    --       .readdata
			m_write         => sd_cont_0_master_write,                       --       .write
			m_writedata     => sd_cont_0_master_writedata,                   --       .writedata
			m_waitrequest_n => sd_cont_0_master_inv,                         --       .waitrequest_n
			sd_clk          => sd_sd_clk,                                    --     sd.sd_clk
			sd_cmd          => sd_sd_cmd,                                    --       .sd_cmd
			sd_dat          => sd_sd_dat,                                    --       .sd_dat
			sd_pll_clk      => clk_50_clk                                    -- sd_clk.clk
		);

	sram : component HW_QSYS_sram
		generic map (
			TCM_ADDRESS_W                  => 19,
			TCM_DATA_W                     => 16,
			TCM_BYTEENABLE_W               => 2,
			TCM_READ_WAIT                  => 10,
			TCM_WRITE_WAIT                 => 10,
			TCM_SETUP_WAIT                 => 10,
			TCM_DATA_HOLD                  => 10,
			TCM_TURNAROUND_TIME            => 2,
			TCM_TIMING_UNITS               => 0,
			TCM_READLATENCY                => 2,
			TCM_SYMBOLS_PER_WORD           => 2,
			USE_READDATA                   => 1,
			USE_WRITEDATA                  => 1,
			USE_READ                       => 0,
			USE_WRITE                      => 1,
			USE_BYTEENABLE                 => 1,
			USE_CHIPSELECT                 => 1,
			USE_LOCK                       => 0,
			USE_ADDRESS                    => 1,
			USE_WAITREQUEST                => 0,
			USE_WRITEBYTEENABLE            => 0,
			USE_OUTPUTENABLE               => 1,
			USE_RESETREQUEST               => 0,
			USE_IRQ                        => 0,
			USE_RESET_OUTPUT               => 0,
			ACTIVE_LOW_READ                => 0,
			ACTIVE_LOW_LOCK                => 0,
			ACTIVE_LOW_WRITE               => 1,
			ACTIVE_LOW_CHIPSELECT          => 1,
			ACTIVE_LOW_BYTEENABLE          => 1,
			ACTIVE_LOW_OUTPUTENABLE        => 1,
			ACTIVE_LOW_WRITEBYTEENABLE     => 0,
			ACTIVE_LOW_WAITREQUEST         => 0,
			ACTIVE_LOW_BEGINTRANSFER       => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0
		)
		port map (
			clk_clk                => clk_125_clk,                              --   clk.clk
			reset_reset            => rst_controller_004_reset_out_reset,       -- reset.reset
			uas_address            => mm_interconnect_0_sram_uas_address,       --   uas.address
			uas_burstcount         => mm_interconnect_0_sram_uas_burstcount,    --      .burstcount
			uas_read               => mm_interconnect_0_sram_uas_read,          --      .read
			uas_write              => mm_interconnect_0_sram_uas_write,         --      .write
			uas_waitrequest        => mm_interconnect_0_sram_uas_waitrequest,   --      .waitrequest
			uas_readdatavalid      => mm_interconnect_0_sram_uas_readdatavalid, --      .readdatavalid
			uas_byteenable         => mm_interconnect_0_sram_uas_byteenable,    --      .byteenable
			uas_readdata           => mm_interconnect_0_sram_uas_readdata,      --      .readdata
			uas_writedata          => mm_interconnect_0_sram_uas_writedata,     --      .writedata
			uas_lock               => mm_interconnect_0_sram_uas_lock,          --      .lock
			uas_debugaccess        => mm_interconnect_0_sram_uas_debugaccess,   --      .debugaccess
			tcm_write_n_out        => sram_tcm_write_n_out,                     --   tcm.write_n_out
			tcm_chipselect_n_out   => sram_tcm_chipselect_n_out,                --      .chipselect_n_out
			tcm_outputenable_n_out => sram_tcm_outputenable_n_out,              --      .outputenable_n_out
			tcm_request            => sram_tcm_request,                         --      .request
			tcm_grant              => sram_tcm_grant,                           --      .grant
			tcm_address_out        => sram_tcm_address_out,                     --      .address_out
			tcm_byteenable_n_out   => sram_tcm_byteenable_n_out,                --      .byteenable_n_out
			tcm_data_out           => sram_tcm_data_out,                        --      .data_out
			tcm_data_outen         => sram_tcm_data_outen,                      --      .data_outen
			tcm_data_in            => sram_tcm_data_in                          --      .data_in
		);

	sram_bridge : component HW_QSYS_sram_bridge
		port map (
			clk                             => clk_125_clk,                                     --   clk.clk
			reset                           => rst_controller_004_reset_out_reset,              -- reset.reset
			request                         => sram_sharer_tcm_request,                         --   tcs.request
			grant                           => sram_sharer_tcm_grant,                           --      .grant
			tcs_sram_tcm_data_out           => sram_sharer_tcm_sram_tcm_data_out_out,           --      .sram_tcm_data_out_out
			tcs_sram_tcm_data_outen         => sram_sharer_tcm_sram_tcm_data_out_outen,         --      .sram_tcm_data_out_outen
			tcs_sram_tcm_data_in            => sram_sharer_tcm_sram_tcm_data_out_in,            --      .sram_tcm_data_out_in
			tcs_sram_tcm_address_out        => sram_sharer_tcm_sram_tcm_address_out_out,        --      .sram_tcm_address_out_out
			tcs_sram_tcm_outputenable_n_out => sram_sharer_tcm_sram_tcm_outputenable_n_out_out, --      .sram_tcm_outputenable_n_out_out
			tcs_sram_tcm_chipselect_n_out   => sram_sharer_tcm_sram_tcm_chipselect_n_out_out,   --      .sram_tcm_chipselect_n_out_out
			tcs_sram_tcm_byteenable_n_out   => sram_sharer_tcm_sram_tcm_byteenable_n_out_out,   --      .sram_tcm_byteenable_n_out_out
			tcs_sram_tcm_write_n_out        => sram_sharer_tcm_sram_tcm_write_n_out_out,        --      .sram_tcm_write_n_out_out
			sram_tcm_data_out               => sram_bridge_out_sram_tcm_data_out,               --   out.sram_tcm_data_out
			sram_tcm_address_out            => sram_bridge_out_sram_tcm_address_out,            --      .sram_tcm_address_out
			sram_tcm_outputenable_n_out     => sram_bridge_out_sram_tcm_outputenable_n_out,     --      .sram_tcm_outputenable_n_out
			sram_tcm_chipselect_n_out       => sram_bridge_out_sram_tcm_chipselect_n_out,       --      .sram_tcm_chipselect_n_out
			sram_tcm_byteenable_n_out       => sram_bridge_out_sram_tcm_byteenable_n_out,       --      .sram_tcm_byteenable_n_out
			sram_tcm_write_n_out            => sram_bridge_out_sram_tcm_write_n_out             --      .sram_tcm_write_n_out
		);

	sram_sharer : component HW_QSYS_sram_sharer
		port map (
			clk_clk                     => clk_125_clk,                                     --   clk.clk
			reset_reset                 => rst_controller_004_reset_out_reset,              -- reset.reset
			request                     => sram_sharer_tcm_request,                         --   tcm.request
			grant                       => sram_sharer_tcm_grant,                           --      .grant
			sram_tcm_address_out        => sram_sharer_tcm_sram_tcm_address_out_out,        --      .sram_tcm_address_out_out
			sram_tcm_byteenable_n_out   => sram_sharer_tcm_sram_tcm_byteenable_n_out_out,   --      .sram_tcm_byteenable_n_out_out
			sram_tcm_outputenable_n_out => sram_sharer_tcm_sram_tcm_outputenable_n_out_out, --      .sram_tcm_outputenable_n_out_out
			sram_tcm_write_n_out        => sram_sharer_tcm_sram_tcm_write_n_out_out,        --      .sram_tcm_write_n_out_out
			sram_tcm_data_out           => sram_sharer_tcm_sram_tcm_data_out_out,           --      .sram_tcm_data_out_out
			sram_tcm_data_in            => sram_sharer_tcm_sram_tcm_data_out_in,            --      .sram_tcm_data_out_in
			sram_tcm_data_outen         => sram_sharer_tcm_sram_tcm_data_out_outen,         --      .sram_tcm_data_out_outen
			sram_tcm_chipselect_n_out   => sram_sharer_tcm_sram_tcm_chipselect_n_out_out,   --      .sram_tcm_chipselect_n_out_out
			tcs0_request                => sram_tcm_request,                                --  tcs0.request
			tcs0_grant                  => sram_tcm_grant,                                  --      .grant
			tcs0_address_out            => sram_tcm_address_out,                            --      .address_out
			tcs0_byteenable_n_out       => sram_tcm_byteenable_n_out,                       --      .byteenable_n_out
			tcs0_outputenable_n_out(0)  => sram_tcm_outputenable_n_out,                     --      .outputenable_n_out
			tcs0_write_n_out(0)         => sram_tcm_write_n_out,                            --      .write_n_out
			tcs0_data_out               => sram_tcm_data_out,                               --      .data_out
			tcs0_data_in                => sram_tcm_data_in,                                --      .data_in
			tcs0_data_outen             => sram_tcm_data_outen,                             --      .data_outen
			tcs0_chipselect_n_out(0)    => sram_tcm_chipselect_n_out                        --      .chipselect_n_out
		);

	sysid : component HW_QSYS_sysid
		port map (
			clock    => clk_125_clk,                                      --           clk.clk
			reset_n  => rst_controller_004_reset_out_reset_ports_inv,     --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	timer_0 : component HW_QSYS_timer_0
		port map (
			clk        => clk_125_clk,                                  --   clk.clk
			reset_n    => rst_controller_004_reset_out_reset_ports_inv, -- reset.reset_n
			address    => mm_interconnect_0_timer_0_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_0_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_0_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_0_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_0_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver5_irq                      --   irq.irq
		);

	timer_1 : component HW_QSYS_timer_1
		port map (
			clk        => clk_125_clk,                                  --   clk.clk
			reset_n    => rst_controller_004_reset_out_reset_ports_inv, -- reset.reset_n
			address    => mm_interconnect_0_timer_1_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_1_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_1_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_1_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_1_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver8_irq                      --   irq.irq
		);

	twod_idct_st_hw_0 : component twod_idct_st_hw
		port map (
			CLOCK     => clk_125_clk,                        -- clock.clk
			DATAOUT   => twod_idct_st_hw_0_dst_data,         --   dst.data
			dst_ready => twod_idct_st_hw_0_dst_ready,        --      .ready
			dst_valid => twod_idct_st_hw_0_dst_valid,        --      .valid
			reset     => rst_controller_004_reset_out_reset, -- reset.reset
			DATAIN    => read_dma_0_st_source_data,          --   src.data
			src_ready => read_dma_0_st_source_ready,         --      .ready
			src_valid => read_dma_0_st_source_valid          --      .valid
		);

	video : component altera_avalon_video_sync_generator
		generic map (
			DATA_STREAM_BIT_WIDTH => 24,
			BEATS_PER_PIXEL       => 1,
			NUM_COLUMNS           => 640,
			NUM_ROWS              => 480,
			H_BLANK_PIXELS        => 128,
			H_FRONT_PORCH_PIXELS  => 24,
			H_SYNC_PULSE_PIXELS   => 32,
			H_SYNC_PULSE_POLARITY => 0,
			V_BLANK_LINES         => 45,
			V_FRONT_PORCH_LINES   => 10,
			V_SYNC_PULSE_LINES    => 3,
			V_SYNC_PULSE_POLARITY => 0,
			TOTAL_HSCAN_PIXELS    => 768,
			TOTAL_VSCAN_LINES     => 525
		)
		port map (
			clk     => video_pll_outclk0_clk,                    --       clk.clk
			reset_n => rst_controller_reset_out_reset_ports_inv, -- clk_reset.reset_n
			ready   => pixel_con_out_ready,                      --        in.ready
			valid   => pixel_con_out_valid,                      --          .valid
			data    => pixel_con_out_data,                       --          .data
			eop     => pixel_con_out_endofpacket,                --          .endofpacket
			sop     => pixel_con_out_startofpacket,              --          .startofpacket
			empty   => pixel_con_out_empty,                      --          .empty
			RGB_OUT => video_RGB_OUT,                            --      sync.export
			HD      => video_HD,                                 --          .export
			VD      => video_VD,                                 --          .export
			DEN     => video_DEN                                 --          .export
		);

	video_dma : component HW_QSYS_video_dma
		port map (
			mm_read_address              => video_dma_mm_read_address,                                --          mm_read.address
			mm_read_read                 => video_dma_mm_read_read,                                   --                 .read
			mm_read_byteenable           => video_dma_mm_read_byteenable,                             --                 .byteenable
			mm_read_readdata             => video_dma_mm_read_readdata,                               --                 .readdata
			mm_read_waitrequest          => video_dma_mm_read_waitrequest,                            --                 .waitrequest
			mm_read_readdatavalid        => video_dma_mm_read_readdatavalid,                          --                 .readdatavalid
			mm_read_burstcount           => video_dma_mm_read_burstcount,                             --                 .burstcount
			clock_clk                    => clk_125_clk,                                              --            clock.clk
			reset_n_reset_n              => rst_controller_004_reset_out_reset_ports_inv,             --          reset_n.reset_n
			csr_writedata                => mm_interconnect_0_video_dma_csr_writedata,                --              csr.writedata
			csr_write                    => mm_interconnect_0_video_dma_csr_write,                    --                 .write
			csr_byteenable               => mm_interconnect_0_video_dma_csr_byteenable,               --                 .byteenable
			csr_readdata                 => mm_interconnect_0_video_dma_csr_readdata,                 --                 .readdata
			csr_read                     => mm_interconnect_0_video_dma_csr_read,                     --                 .read
			csr_address                  => mm_interconnect_0_video_dma_csr_address,                  --                 .address
			descriptor_slave_write       => mm_interconnect_0_video_dma_descriptor_slave_write,       -- descriptor_slave.write
			descriptor_slave_waitrequest => mm_interconnect_0_video_dma_descriptor_slave_waitrequest, --                 .waitrequest
			descriptor_slave_writedata   => mm_interconnect_0_video_dma_descriptor_slave_writedata,   --                 .writedata
			descriptor_slave_byteenable  => mm_interconnect_0_video_dma_descriptor_slave_byteenable,  --                 .byteenable
			csr_irq_irq                  => irq_mapper_receiver0_irq,                                 --          csr_irq.irq
			st_source_data               => video_dma_st_source_data,                                 --        st_source.data
			st_source_valid              => video_dma_st_source_valid,                                --                 .valid
			st_source_ready              => video_dma_st_source_ready,                                --                 .ready
			st_source_startofpacket      => video_dma_st_source_startofpacket,                        --                 .startofpacket
			st_source_endofpacket        => video_dma_st_source_endofpacket,                          --                 .endofpacket
			st_source_empty              => video_dma_st_source_empty                                 --                 .empty
		);

	video_fifo : component HW_QSYS_video_fifo
		port map (
			wrclock                       => clk_125_clk,                                  --    clk_in.clk
			wrreset_n                     => rst_controller_004_reset_out_reset_ports_inv, --  reset_in.reset_n
			rdclock                       => video_pll_outclk0_clk,                        --   clk_out.clk
			rdreset_n                     => rst_controller_reset_out_reset_ports_inv,     -- reset_out.reset_n
			avalonst_sink_valid           => avalon_st_adapter_001_out_0_valid,            --        in.valid
			avalonst_sink_data            => avalon_st_adapter_001_out_0_data,             --          .data
			avalonst_sink_startofpacket   => avalon_st_adapter_001_out_0_startofpacket,    --          .startofpacket
			avalonst_sink_endofpacket     => avalon_st_adapter_001_out_0_endofpacket,      --          .endofpacket
			avalonst_sink_empty           => avalon_st_adapter_001_out_0_empty,            --          .empty
			avalonst_sink_ready           => avalon_st_adapter_001_out_0_ready,            --          .ready
			avalonst_source_valid         => video_fifo_out_valid,                         --       out.valid
			avalonst_source_data          => video_fifo_out_data,                          --          .data
			avalonst_source_startofpacket => video_fifo_out_startofpacket,                 --          .startofpacket
			avalonst_source_endofpacket   => video_fifo_out_endofpacket,                   --          .endofpacket
			avalonst_source_empty         => video_fifo_out_empty,                         --          .empty
			avalonst_source_ready         => video_fifo_out_ready                          --          .ready
		);

	video_pll : component HW_QSYS_video_pll
		port map (
			refclk   => clk_50_clk,                         --  refclk.clk
			rst      => reset_controller_0_reset_out_reset, --   reset.reset
			outclk_0 => video_pll_outclk0_clk,              -- outclk0.clk
			locked   => open                                -- (terminated)
		);

	write_dma_0 : component HW_QSYS_write_dma_0
		port map (
			mm_write_address             => write_dma_0_mm_write_address,                               --         mm_write.address
			mm_write_write               => write_dma_0_mm_write_write,                                 --                 .write
			mm_write_byteenable          => write_dma_0_mm_write_byteenable,                            --                 .byteenable
			mm_write_writedata           => write_dma_0_mm_write_writedata,                             --                 .writedata
			mm_write_waitrequest         => write_dma_0_mm_write_waitrequest,                           --                 .waitrequest
			mm_write_burstcount          => write_dma_0_mm_write_burstcount,                            --                 .burstcount
			clock_clk                    => clk_125_clk,                                                --            clock.clk
			reset_n_reset_n              => rst_controller_004_reset_out_reset_ports_inv,               --          reset_n.reset_n
			csr_writedata                => mm_interconnect_0_write_dma_0_csr_writedata,                --              csr.writedata
			csr_write                    => mm_interconnect_0_write_dma_0_csr_write,                    --                 .write
			csr_byteenable               => mm_interconnect_0_write_dma_0_csr_byteenable,               --                 .byteenable
			csr_readdata                 => mm_interconnect_0_write_dma_0_csr_readdata,                 --                 .readdata
			csr_read                     => mm_interconnect_0_write_dma_0_csr_read,                     --                 .read
			csr_address                  => mm_interconnect_0_write_dma_0_csr_address,                  --                 .address
			descriptor_slave_write       => mm_interconnect_0_write_dma_0_descriptor_slave_write,       -- descriptor_slave.write
			descriptor_slave_waitrequest => mm_interconnect_0_write_dma_0_descriptor_slave_waitrequest, --                 .waitrequest
			descriptor_slave_writedata   => mm_interconnect_0_write_dma_0_descriptor_slave_writedata,   --                 .writedata
			descriptor_slave_byteenable  => mm_interconnect_0_write_dma_0_descriptor_slave_byteenable,  --                 .byteenable
			csr_irq_irq                  => irq_mapper_receiver1_irq,                                   --          csr_irq.irq
			st_sink_data                 => twod_idct_st_hw_0_dst_data,                                 --          st_sink.data
			st_sink_valid                => twod_idct_st_hw_0_dst_valid,                                --                 .valid
			st_sink_ready                => twod_idct_st_hw_0_dst_ready                                 --                 .ready
		);

	mm_interconnect_0 : component HW_QSYS_mm_interconnect_0
		port map (
			clk_125_clk_clk                                     => clk_125_clk,                                                    --                                   clk_125_clk.clk
			clk_50_out_clk_clk                                  => clk_50_clk,                                                     --                                clk_50_out_clk.clk
			cpu_0_reset_reset_bridge_in_reset_reset             => rst_controller_001_reset_out_reset,                             --             cpu_0_reset_reset_bridge_in_reset.reset
			cpu_1_reset_reset_bridge_in_reset_reset             => rst_controller_002_reset_out_reset,                             --             cpu_1_reset_reset_bridge_in_reset.reset
			cpu_2_reset_reset_bridge_in_reset_reset             => rst_controller_003_reset_out_reset,                             --             cpu_2_reset_reset_bridge_in_reset.reset
			lpddr2_mp_cmd_reset_n_0_reset_bridge_in_reset_reset => rst_controller_004_reset_out_reset,                             -- lpddr2_mp_cmd_reset_n_0_reset_bridge_in_reset.reset
			mailbox_simple_1_rst_n_reset_bridge_in_reset_reset  => rst_controller_004_reset_out_reset,                             --  mailbox_simple_1_rst_n_reset_bridge_in_reset.reset
			sd_cont_0_reset_reset_bridge_in_reset_reset         => rst_controller_005_reset_out_reset,                             --         sd_cont_0_reset_reset_bridge_in_reset.reset
			cpu_0_data_master_address                           => cpu_0_data_master_address,                                      --                             cpu_0_data_master.address
			cpu_0_data_master_waitrequest                       => cpu_0_data_master_waitrequest,                                  --                                              .waitrequest
			cpu_0_data_master_burstcount                        => cpu_0_data_master_burstcount,                                   --                                              .burstcount
			cpu_0_data_master_byteenable                        => cpu_0_data_master_byteenable,                                   --                                              .byteenable
			cpu_0_data_master_read                              => cpu_0_data_master_read,                                         --                                              .read
			cpu_0_data_master_readdata                          => cpu_0_data_master_readdata,                                     --                                              .readdata
			cpu_0_data_master_readdatavalid                     => cpu_0_data_master_readdatavalid,                                --                                              .readdatavalid
			cpu_0_data_master_write                             => cpu_0_data_master_write,                                        --                                              .write
			cpu_0_data_master_writedata                         => cpu_0_data_master_writedata,                                    --                                              .writedata
			cpu_0_data_master_debugaccess                       => cpu_0_data_master_debugaccess,                                  --                                              .debugaccess
			cpu_0_instruction_master_address                    => cpu_0_instruction_master_address,                               --                      cpu_0_instruction_master.address
			cpu_0_instruction_master_waitrequest                => cpu_0_instruction_master_waitrequest,                           --                                              .waitrequest
			cpu_0_instruction_master_read                       => cpu_0_instruction_master_read,                                  --                                              .read
			cpu_0_instruction_master_readdata                   => cpu_0_instruction_master_readdata,                              --                                              .readdata
			cpu_0_instruction_master_readdatavalid              => cpu_0_instruction_master_readdatavalid,                         --                                              .readdatavalid
			cpu_1_data_master_address                           => cpu_1_data_master_address,                                      --                             cpu_1_data_master.address
			cpu_1_data_master_waitrequest                       => cpu_1_data_master_waitrequest,                                  --                                              .waitrequest
			cpu_1_data_master_burstcount                        => cpu_1_data_master_burstcount,                                   --                                              .burstcount
			cpu_1_data_master_byteenable                        => cpu_1_data_master_byteenable,                                   --                                              .byteenable
			cpu_1_data_master_read                              => cpu_1_data_master_read,                                         --                                              .read
			cpu_1_data_master_readdata                          => cpu_1_data_master_readdata,                                     --                                              .readdata
			cpu_1_data_master_readdatavalid                     => cpu_1_data_master_readdatavalid,                                --                                              .readdatavalid
			cpu_1_data_master_write                             => cpu_1_data_master_write,                                        --                                              .write
			cpu_1_data_master_writedata                         => cpu_1_data_master_writedata,                                    --                                              .writedata
			cpu_1_data_master_debugaccess                       => cpu_1_data_master_debugaccess,                                  --                                              .debugaccess
			cpu_1_instruction_master_address                    => cpu_1_instruction_master_address,                               --                      cpu_1_instruction_master.address
			cpu_1_instruction_master_waitrequest                => cpu_1_instruction_master_waitrequest,                           --                                              .waitrequest
			cpu_1_instruction_master_read                       => cpu_1_instruction_master_read,                                  --                                              .read
			cpu_1_instruction_master_readdata                   => cpu_1_instruction_master_readdata,                              --                                              .readdata
			cpu_1_instruction_master_readdatavalid              => cpu_1_instruction_master_readdatavalid,                         --                                              .readdatavalid
			cpu_2_data_master_address                           => cpu_2_data_master_address,                                      --                             cpu_2_data_master.address
			cpu_2_data_master_waitrequest                       => cpu_2_data_master_waitrequest,                                  --                                              .waitrequest
			cpu_2_data_master_burstcount                        => cpu_2_data_master_burstcount,                                   --                                              .burstcount
			cpu_2_data_master_byteenable                        => cpu_2_data_master_byteenable,                                   --                                              .byteenable
			cpu_2_data_master_read                              => cpu_2_data_master_read,                                         --                                              .read
			cpu_2_data_master_readdata                          => cpu_2_data_master_readdata,                                     --                                              .readdata
			cpu_2_data_master_readdatavalid                     => cpu_2_data_master_readdatavalid,                                --                                              .readdatavalid
			cpu_2_data_master_write                             => cpu_2_data_master_write,                                        --                                              .write
			cpu_2_data_master_writedata                         => cpu_2_data_master_writedata,                                    --                                              .writedata
			cpu_2_data_master_debugaccess                       => cpu_2_data_master_debugaccess,                                  --                                              .debugaccess
			cpu_2_instruction_master_address                    => cpu_2_instruction_master_address,                               --                      cpu_2_instruction_master.address
			cpu_2_instruction_master_waitrequest                => cpu_2_instruction_master_waitrequest,                           --                                              .waitrequest
			cpu_2_instruction_master_read                       => cpu_2_instruction_master_read,                                  --                                              .read
			cpu_2_instruction_master_readdata                   => cpu_2_instruction_master_readdata,                              --                                              .readdata
			cpu_2_instruction_master_readdatavalid              => cpu_2_instruction_master_readdatavalid,                         --                                              .readdatavalid
			sd_cont_0_master_address                            => sd_cont_0_master_address,                                       --                              sd_cont_0_master.address
			sd_cont_0_master_waitrequest                        => mm_interconnect_0_sd_cont_0_master_waitrequest,                 --                                              .waitrequest
			sd_cont_0_master_read                               => sd_cont_0_master_read,                                          --                                              .read
			sd_cont_0_master_readdata                           => sd_cont_0_master_readdata,                                      --                                              .readdata
			sd_cont_0_master_write                              => sd_cont_0_master_write,                                         --                                              .write
			sd_cont_0_master_writedata                          => sd_cont_0_master_writedata,                                     --                                              .writedata
			cpu_0_debug_mem_slave_address                       => mm_interconnect_0_cpu_0_debug_mem_slave_address,                --                         cpu_0_debug_mem_slave.address
			cpu_0_debug_mem_slave_write                         => mm_interconnect_0_cpu_0_debug_mem_slave_write,                  --                                              .write
			cpu_0_debug_mem_slave_read                          => mm_interconnect_0_cpu_0_debug_mem_slave_read,                   --                                              .read
			cpu_0_debug_mem_slave_readdata                      => mm_interconnect_0_cpu_0_debug_mem_slave_readdata,               --                                              .readdata
			cpu_0_debug_mem_slave_writedata                     => mm_interconnect_0_cpu_0_debug_mem_slave_writedata,              --                                              .writedata
			cpu_0_debug_mem_slave_byteenable                    => mm_interconnect_0_cpu_0_debug_mem_slave_byteenable,             --                                              .byteenable
			cpu_0_debug_mem_slave_waitrequest                   => mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest,            --                                              .waitrequest
			cpu_0_debug_mem_slave_debugaccess                   => mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess,            --                                              .debugaccess
			cpu_1_debug_mem_slave_address                       => mm_interconnect_0_cpu_1_debug_mem_slave_address,                --                         cpu_1_debug_mem_slave.address
			cpu_1_debug_mem_slave_write                         => mm_interconnect_0_cpu_1_debug_mem_slave_write,                  --                                              .write
			cpu_1_debug_mem_slave_read                          => mm_interconnect_0_cpu_1_debug_mem_slave_read,                   --                                              .read
			cpu_1_debug_mem_slave_readdata                      => mm_interconnect_0_cpu_1_debug_mem_slave_readdata,               --                                              .readdata
			cpu_1_debug_mem_slave_writedata                     => mm_interconnect_0_cpu_1_debug_mem_slave_writedata,              --                                              .writedata
			cpu_1_debug_mem_slave_byteenable                    => mm_interconnect_0_cpu_1_debug_mem_slave_byteenable,             --                                              .byteenable
			cpu_1_debug_mem_slave_waitrequest                   => mm_interconnect_0_cpu_1_debug_mem_slave_waitrequest,            --                                              .waitrequest
			cpu_1_debug_mem_slave_debugaccess                   => mm_interconnect_0_cpu_1_debug_mem_slave_debugaccess,            --                                              .debugaccess
			cpu_2_debug_mem_slave_address                       => mm_interconnect_0_cpu_2_debug_mem_slave_address,                --                         cpu_2_debug_mem_slave.address
			cpu_2_debug_mem_slave_write                         => mm_interconnect_0_cpu_2_debug_mem_slave_write,                  --                                              .write
			cpu_2_debug_mem_slave_read                          => mm_interconnect_0_cpu_2_debug_mem_slave_read,                   --                                              .read
			cpu_2_debug_mem_slave_readdata                      => mm_interconnect_0_cpu_2_debug_mem_slave_readdata,               --                                              .readdata
			cpu_2_debug_mem_slave_writedata                     => mm_interconnect_0_cpu_2_debug_mem_slave_writedata,              --                                              .writedata
			cpu_2_debug_mem_slave_byteenable                    => mm_interconnect_0_cpu_2_debug_mem_slave_byteenable,             --                                              .byteenable
			cpu_2_debug_mem_slave_waitrequest                   => mm_interconnect_0_cpu_2_debug_mem_slave_waitrequest,            --                                              .waitrequest
			cpu_2_debug_mem_slave_debugaccess                   => mm_interconnect_0_cpu_2_debug_mem_slave_debugaccess,            --                                              .debugaccess
			i2c_scl_s1_address                                  => mm_interconnect_0_i2c_scl_s1_address,                           --                                    i2c_scl_s1.address
			i2c_scl_s1_write                                    => mm_interconnect_0_i2c_scl_s1_write,                             --                                              .write
			i2c_scl_s1_readdata                                 => mm_interconnect_0_i2c_scl_s1_readdata,                          --                                              .readdata
			i2c_scl_s1_writedata                                => mm_interconnect_0_i2c_scl_s1_writedata,                         --                                              .writedata
			i2c_scl_s1_chipselect                               => mm_interconnect_0_i2c_scl_s1_chipselect,                        --                                              .chipselect
			i2c_sda_s1_address                                  => mm_interconnect_0_i2c_sda_s1_address,                           --                                    i2c_sda_s1.address
			i2c_sda_s1_write                                    => mm_interconnect_0_i2c_sda_s1_write,                             --                                              .write
			i2c_sda_s1_readdata                                 => mm_interconnect_0_i2c_sda_s1_readdata,                          --                                              .readdata
			i2c_sda_s1_writedata                                => mm_interconnect_0_i2c_sda_s1_writedata,                         --                                              .writedata
			i2c_sda_s1_chipselect                               => mm_interconnect_0_i2c_sda_s1_chipselect,                        --                                              .chipselect
			jtag_uart_0_avalon_jtag_slave_address               => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,        --                 jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write                 => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,          --                                              .write
			jtag_uart_0_avalon_jtag_slave_read                  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,           --                                              .read
			jtag_uart_0_avalon_jtag_slave_readdata              => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,       --                                              .readdata
			jtag_uart_0_avalon_jtag_slave_writedata             => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,      --                                              .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest           => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,    --                                              .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect            => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,     --                                              .chipselect
			jtag_uart_1_avalon_jtag_slave_address               => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_address,        --                 jtag_uart_1_avalon_jtag_slave.address
			jtag_uart_1_avalon_jtag_slave_write                 => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write,          --                                              .write
			jtag_uart_1_avalon_jtag_slave_read                  => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read,           --                                              .read
			jtag_uart_1_avalon_jtag_slave_readdata              => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_readdata,       --                                              .readdata
			jtag_uart_1_avalon_jtag_slave_writedata             => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_writedata,      --                                              .writedata
			jtag_uart_1_avalon_jtag_slave_waitrequest           => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_waitrequest,    --                                              .waitrequest
			jtag_uart_1_avalon_jtag_slave_chipselect            => mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_chipselect,     --                                              .chipselect
			jtag_uart_2_avalon_jtag_slave_address               => mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_address,        --                 jtag_uart_2_avalon_jtag_slave.address
			jtag_uart_2_avalon_jtag_slave_write                 => mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_write,          --                                              .write
			jtag_uart_2_avalon_jtag_slave_read                  => mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_read,           --                                              .read
			jtag_uart_2_avalon_jtag_slave_readdata              => mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_readdata,       --                                              .readdata
			jtag_uart_2_avalon_jtag_slave_writedata             => mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_writedata,      --                                              .writedata
			jtag_uart_2_avalon_jtag_slave_waitrequest           => mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_waitrequest,    --                                              .waitrequest
			jtag_uart_2_avalon_jtag_slave_chipselect            => mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_chipselect,     --                                              .chipselect
			key_s1_address                                      => mm_interconnect_0_key_s1_address,                               --                                        key_s1.address
			key_s1_write                                        => mm_interconnect_0_key_s1_write,                                 --                                              .write
			key_s1_readdata                                     => mm_interconnect_0_key_s1_readdata,                              --                                              .readdata
			key_s1_writedata                                    => mm_interconnect_0_key_s1_writedata,                             --                                              .writedata
			key_s1_chipselect                                   => mm_interconnect_0_key_s1_chipselect,                            --                                              .chipselect
			ledg_s1_address                                     => mm_interconnect_0_ledg_s1_address,                              --                                       ledg_s1.address
			ledg_s1_write                                       => mm_interconnect_0_ledg_s1_write,                                --                                              .write
			ledg_s1_readdata                                    => mm_interconnect_0_ledg_s1_readdata,                             --                                              .readdata
			ledg_s1_writedata                                   => mm_interconnect_0_ledg_s1_writedata,                            --                                              .writedata
			ledg_s1_chipselect                                  => mm_interconnect_0_ledg_s1_chipselect,                           --                                              .chipselect
			ledr_s1_address                                     => mm_interconnect_0_ledr_s1_address,                              --                                       ledr_s1.address
			ledr_s1_write                                       => mm_interconnect_0_ledr_s1_write,                                --                                              .write
			ledr_s1_readdata                                    => mm_interconnect_0_ledr_s1_readdata,                             --                                              .readdata
			ledr_s1_writedata                                   => mm_interconnect_0_ledr_s1_writedata,                            --                                              .writedata
			ledr_s1_chipselect                                  => mm_interconnect_0_ledr_s1_chipselect,                           --                                              .chipselect
			lpddr2_avl_0_address                                => mm_interconnect_0_lpddr2_avl_0_address,                         --                                  lpddr2_avl_0.address
			lpddr2_avl_0_write                                  => mm_interconnect_0_lpddr2_avl_0_write,                           --                                              .write
			lpddr2_avl_0_read                                   => mm_interconnect_0_lpddr2_avl_0_read,                            --                                              .read
			lpddr2_avl_0_readdata                               => mm_interconnect_0_lpddr2_avl_0_readdata,                        --                                              .readdata
			lpddr2_avl_0_writedata                              => mm_interconnect_0_lpddr2_avl_0_writedata,                       --                                              .writedata
			lpddr2_avl_0_beginbursttransfer                     => mm_interconnect_0_lpddr2_avl_0_beginbursttransfer,              --                                              .beginbursttransfer
			lpddr2_avl_0_burstcount                             => mm_interconnect_0_lpddr2_avl_0_burstcount,                      --                                              .burstcount
			lpddr2_avl_0_byteenable                             => mm_interconnect_0_lpddr2_avl_0_byteenable,                      --                                              .byteenable
			lpddr2_avl_0_readdatavalid                          => mm_interconnect_0_lpddr2_avl_0_readdatavalid,                   --                                              .readdatavalid
			lpddr2_avl_0_waitrequest                            => mm_interconnect_0_lpddr2_avl_0_inv,                             --                                              .waitrequest
			mailbox_simple_0_avmm_msg_receiver_address          => mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_address,   --            mailbox_simple_0_avmm_msg_receiver.address
			mailbox_simple_0_avmm_msg_receiver_write            => mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_write,     --                                              .write
			mailbox_simple_0_avmm_msg_receiver_read             => mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_read,      --                                              .read
			mailbox_simple_0_avmm_msg_receiver_readdata         => mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_readdata,  --                                              .readdata
			mailbox_simple_0_avmm_msg_receiver_writedata        => mm_interconnect_0_mailbox_simple_0_avmm_msg_receiver_writedata, --                                              .writedata
			mailbox_simple_0_avmm_msg_sender_address            => mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_address,     --              mailbox_simple_0_avmm_msg_sender.address
			mailbox_simple_0_avmm_msg_sender_write              => mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_write,       --                                              .write
			mailbox_simple_0_avmm_msg_sender_read               => mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_read,        --                                              .read
			mailbox_simple_0_avmm_msg_sender_readdata           => mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_readdata,    --                                              .readdata
			mailbox_simple_0_avmm_msg_sender_writedata          => mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_writedata,   --                                              .writedata
			mailbox_simple_0_avmm_msg_sender_waitrequest        => mm_interconnect_0_mailbox_simple_0_avmm_msg_sender_waitrequest, --                                              .waitrequest
			mailbox_simple_1_avmm_msg_receiver_address          => mm_interconnect_0_mailbox_simple_1_avmm_msg_receiver_address,   --            mailbox_simple_1_avmm_msg_receiver.address
			mailbox_simple_1_avmm_msg_receiver_write            => mm_interconnect_0_mailbox_simple_1_avmm_msg_receiver_write,     --                                              .write
			mailbox_simple_1_avmm_msg_receiver_read             => mm_interconnect_0_mailbox_simple_1_avmm_msg_receiver_read,      --                                              .read
			mailbox_simple_1_avmm_msg_receiver_readdata         => mm_interconnect_0_mailbox_simple_1_avmm_msg_receiver_readdata,  --                                              .readdata
			mailbox_simple_1_avmm_msg_receiver_writedata        => mm_interconnect_0_mailbox_simple_1_avmm_msg_receiver_writedata, --                                              .writedata
			mailbox_simple_1_avmm_msg_sender_address            => mm_interconnect_0_mailbox_simple_1_avmm_msg_sender_address,     --              mailbox_simple_1_avmm_msg_sender.address
			mailbox_simple_1_avmm_msg_sender_write              => mm_interconnect_0_mailbox_simple_1_avmm_msg_sender_write,       --                                              .write
			mailbox_simple_1_avmm_msg_sender_read               => mm_interconnect_0_mailbox_simple_1_avmm_msg_sender_read,        --                                              .read
			mailbox_simple_1_avmm_msg_sender_readdata           => mm_interconnect_0_mailbox_simple_1_avmm_msg_sender_readdata,    --                                              .readdata
			mailbox_simple_1_avmm_msg_sender_writedata          => mm_interconnect_0_mailbox_simple_1_avmm_msg_sender_writedata,   --                                              .writedata
			mailbox_simple_1_avmm_msg_sender_waitrequest        => mm_interconnect_0_mailbox_simple_1_avmm_msg_sender_waitrequest, --                                              .waitrequest
			mailbox_simple_2_avmm_msg_receiver_address          => mm_interconnect_0_mailbox_simple_2_avmm_msg_receiver_address,   --            mailbox_simple_2_avmm_msg_receiver.address
			mailbox_simple_2_avmm_msg_receiver_write            => mm_interconnect_0_mailbox_simple_2_avmm_msg_receiver_write,     --                                              .write
			mailbox_simple_2_avmm_msg_receiver_read             => mm_interconnect_0_mailbox_simple_2_avmm_msg_receiver_read,      --                                              .read
			mailbox_simple_2_avmm_msg_receiver_readdata         => mm_interconnect_0_mailbox_simple_2_avmm_msg_receiver_readdata,  --                                              .readdata
			mailbox_simple_2_avmm_msg_receiver_writedata        => mm_interconnect_0_mailbox_simple_2_avmm_msg_receiver_writedata, --                                              .writedata
			mailbox_simple_2_avmm_msg_sender_address            => mm_interconnect_0_mailbox_simple_2_avmm_msg_sender_address,     --              mailbox_simple_2_avmm_msg_sender.address
			mailbox_simple_2_avmm_msg_sender_write              => mm_interconnect_0_mailbox_simple_2_avmm_msg_sender_write,       --                                              .write
			mailbox_simple_2_avmm_msg_sender_read               => mm_interconnect_0_mailbox_simple_2_avmm_msg_sender_read,        --                                              .read
			mailbox_simple_2_avmm_msg_sender_readdata           => mm_interconnect_0_mailbox_simple_2_avmm_msg_sender_readdata,    --                                              .readdata
			mailbox_simple_2_avmm_msg_sender_writedata          => mm_interconnect_0_mailbox_simple_2_avmm_msg_sender_writedata,   --                                              .writedata
			mailbox_simple_2_avmm_msg_sender_waitrequest        => mm_interconnect_0_mailbox_simple_2_avmm_msg_sender_waitrequest, --                                              .waitrequest
			mailbox_simple_3_avmm_msg_receiver_address          => mm_interconnect_0_mailbox_simple_3_avmm_msg_receiver_address,   --            mailbox_simple_3_avmm_msg_receiver.address
			mailbox_simple_3_avmm_msg_receiver_write            => mm_interconnect_0_mailbox_simple_3_avmm_msg_receiver_write,     --                                              .write
			mailbox_simple_3_avmm_msg_receiver_read             => mm_interconnect_0_mailbox_simple_3_avmm_msg_receiver_read,      --                                              .read
			mailbox_simple_3_avmm_msg_receiver_readdata         => mm_interconnect_0_mailbox_simple_3_avmm_msg_receiver_readdata,  --                                              .readdata
			mailbox_simple_3_avmm_msg_receiver_writedata        => mm_interconnect_0_mailbox_simple_3_avmm_msg_receiver_writedata, --                                              .writedata
			mailbox_simple_3_avmm_msg_sender_address            => mm_interconnect_0_mailbox_simple_3_avmm_msg_sender_address,     --              mailbox_simple_3_avmm_msg_sender.address
			mailbox_simple_3_avmm_msg_sender_write              => mm_interconnect_0_mailbox_simple_3_avmm_msg_sender_write,       --                                              .write
			mailbox_simple_3_avmm_msg_sender_read               => mm_interconnect_0_mailbox_simple_3_avmm_msg_sender_read,        --                                              .read
			mailbox_simple_3_avmm_msg_sender_readdata           => mm_interconnect_0_mailbox_simple_3_avmm_msg_sender_readdata,    --                                              .readdata
			mailbox_simple_3_avmm_msg_sender_writedata          => mm_interconnect_0_mailbox_simple_3_avmm_msg_sender_writedata,   --                                              .writedata
			mailbox_simple_3_avmm_msg_sender_waitrequest        => mm_interconnect_0_mailbox_simple_3_avmm_msg_sender_waitrequest, --                                              .waitrequest
			read_dma_0_csr_address                              => mm_interconnect_0_read_dma_0_csr_address,                       --                                read_dma_0_csr.address
			read_dma_0_csr_write                                => mm_interconnect_0_read_dma_0_csr_write,                         --                                              .write
			read_dma_0_csr_read                                 => mm_interconnect_0_read_dma_0_csr_read,                          --                                              .read
			read_dma_0_csr_readdata                             => mm_interconnect_0_read_dma_0_csr_readdata,                      --                                              .readdata
			read_dma_0_csr_writedata                            => mm_interconnect_0_read_dma_0_csr_writedata,                     --                                              .writedata
			read_dma_0_csr_byteenable                           => mm_interconnect_0_read_dma_0_csr_byteenable,                    --                                              .byteenable
			read_dma_0_descriptor_slave_write                   => mm_interconnect_0_read_dma_0_descriptor_slave_write,            --                   read_dma_0_descriptor_slave.write
			read_dma_0_descriptor_slave_writedata               => mm_interconnect_0_read_dma_0_descriptor_slave_writedata,        --                                              .writedata
			read_dma_0_descriptor_slave_byteenable              => mm_interconnect_0_read_dma_0_descriptor_slave_byteenable,       --                                              .byteenable
			read_dma_0_descriptor_slave_waitrequest             => mm_interconnect_0_read_dma_0_descriptor_slave_waitrequest,      --                                              .waitrequest
			sd_cont_0_slave_address                             => mm_interconnect_0_sd_cont_0_slave_address,                      --                               sd_cont_0_slave.address
			sd_cont_0_slave_write                               => mm_interconnect_0_sd_cont_0_slave_write,                        --                                              .write
			sd_cont_0_slave_read                                => mm_interconnect_0_sd_cont_0_slave_read,                         --                                              .read
			sd_cont_0_slave_readdata                            => mm_interconnect_0_sd_cont_0_slave_readdata,                     --                                              .readdata
			sd_cont_0_slave_writedata                           => mm_interconnect_0_sd_cont_0_slave_writedata,                    --                                              .writedata
			sd_cont_0_slave_waitrequest                         => mm_interconnect_0_sd_cont_0_slave_inv,                          --                                              .waitrequest
			sd_cont_0_slave_chipselect                          => mm_interconnect_0_sd_cont_0_slave_chipselect,                   --                                              .chipselect
			sram_uas_address                                    => mm_interconnect_0_sram_uas_address,                             --                                      sram_uas.address
			sram_uas_write                                      => mm_interconnect_0_sram_uas_write,                               --                                              .write
			sram_uas_read                                       => mm_interconnect_0_sram_uas_read,                                --                                              .read
			sram_uas_readdata                                   => mm_interconnect_0_sram_uas_readdata,                            --                                              .readdata
			sram_uas_writedata                                  => mm_interconnect_0_sram_uas_writedata,                           --                                              .writedata
			sram_uas_burstcount                                 => mm_interconnect_0_sram_uas_burstcount,                          --                                              .burstcount
			sram_uas_byteenable                                 => mm_interconnect_0_sram_uas_byteenable,                          --                                              .byteenable
			sram_uas_readdatavalid                              => mm_interconnect_0_sram_uas_readdatavalid,                       --                                              .readdatavalid
			sram_uas_waitrequest                                => mm_interconnect_0_sram_uas_waitrequest,                         --                                              .waitrequest
			sram_uas_lock                                       => mm_interconnect_0_sram_uas_lock,                                --                                              .lock
			sram_uas_debugaccess                                => mm_interconnect_0_sram_uas_debugaccess,                         --                                              .debugaccess
			sysid_control_slave_address                         => mm_interconnect_0_sysid_control_slave_address,                  --                           sysid_control_slave.address
			sysid_control_slave_readdata                        => mm_interconnect_0_sysid_control_slave_readdata,                 --                                              .readdata
			timer_0_s1_address                                  => mm_interconnect_0_timer_0_s1_address,                           --                                    timer_0_s1.address
			timer_0_s1_write                                    => mm_interconnect_0_timer_0_s1_write,                             --                                              .write
			timer_0_s1_readdata                                 => mm_interconnect_0_timer_0_s1_readdata,                          --                                              .readdata
			timer_0_s1_writedata                                => mm_interconnect_0_timer_0_s1_writedata,                         --                                              .writedata
			timer_0_s1_chipselect                               => mm_interconnect_0_timer_0_s1_chipselect,                        --                                              .chipselect
			timer_1_s1_address                                  => mm_interconnect_0_timer_1_s1_address,                           --                                    timer_1_s1.address
			timer_1_s1_write                                    => mm_interconnect_0_timer_1_s1_write,                             --                                              .write
			timer_1_s1_readdata                                 => mm_interconnect_0_timer_1_s1_readdata,                          --                                              .readdata
			timer_1_s1_writedata                                => mm_interconnect_0_timer_1_s1_writedata,                         --                                              .writedata
			timer_1_s1_chipselect                               => mm_interconnect_0_timer_1_s1_chipselect,                        --                                              .chipselect
			video_dma_csr_address                               => mm_interconnect_0_video_dma_csr_address,                        --                                 video_dma_csr.address
			video_dma_csr_write                                 => mm_interconnect_0_video_dma_csr_write,                          --                                              .write
			video_dma_csr_read                                  => mm_interconnect_0_video_dma_csr_read,                           --                                              .read
			video_dma_csr_readdata                              => mm_interconnect_0_video_dma_csr_readdata,                       --                                              .readdata
			video_dma_csr_writedata                             => mm_interconnect_0_video_dma_csr_writedata,                      --                                              .writedata
			video_dma_csr_byteenable                            => mm_interconnect_0_video_dma_csr_byteenable,                     --                                              .byteenable
			video_dma_descriptor_slave_write                    => mm_interconnect_0_video_dma_descriptor_slave_write,             --                    video_dma_descriptor_slave.write
			video_dma_descriptor_slave_writedata                => mm_interconnect_0_video_dma_descriptor_slave_writedata,         --                                              .writedata
			video_dma_descriptor_slave_byteenable               => mm_interconnect_0_video_dma_descriptor_slave_byteenable,        --                                              .byteenable
			video_dma_descriptor_slave_waitrequest              => mm_interconnect_0_video_dma_descriptor_slave_waitrequest,       --                                              .waitrequest
			write_dma_0_csr_address                             => mm_interconnect_0_write_dma_0_csr_address,                      --                               write_dma_0_csr.address
			write_dma_0_csr_write                               => mm_interconnect_0_write_dma_0_csr_write,                        --                                              .write
			write_dma_0_csr_read                                => mm_interconnect_0_write_dma_0_csr_read,                         --                                              .read
			write_dma_0_csr_readdata                            => mm_interconnect_0_write_dma_0_csr_readdata,                     --                                              .readdata
			write_dma_0_csr_writedata                           => mm_interconnect_0_write_dma_0_csr_writedata,                    --                                              .writedata
			write_dma_0_csr_byteenable                          => mm_interconnect_0_write_dma_0_csr_byteenable,                   --                                              .byteenable
			write_dma_0_descriptor_slave_write                  => mm_interconnect_0_write_dma_0_descriptor_slave_write,           --                  write_dma_0_descriptor_slave.write
			write_dma_0_descriptor_slave_writedata              => mm_interconnect_0_write_dma_0_descriptor_slave_writedata,       --                                              .writedata
			write_dma_0_descriptor_slave_byteenable             => mm_interconnect_0_write_dma_0_descriptor_slave_byteenable,      --                                              .byteenable
			write_dma_0_descriptor_slave_waitrequest            => mm_interconnect_0_write_dma_0_descriptor_slave_waitrequest      --                                              .waitrequest
		);

	mm_interconnect_1 : component HW_QSYS_mm_interconnect_1
		port map (
			clk_125_clk_clk                                     => clk_125_clk,                                       --                                   clk_125_clk.clk
			lpddr2_mp_cmd_reset_n_1_reset_bridge_in_reset_reset => rst_controller_004_reset_out_reset,                -- lpddr2_mp_cmd_reset_n_1_reset_bridge_in_reset.reset
			video_dma_reset_n_reset_bridge_in_reset_reset       => rst_controller_004_reset_out_reset,                --       video_dma_reset_n_reset_bridge_in_reset.reset
			read_dma_0_mm_read_address                          => read_dma_0_mm_read_address,                        --                            read_dma_0_mm_read.address
			read_dma_0_mm_read_waitrequest                      => read_dma_0_mm_read_waitrequest,                    --                                              .waitrequest
			read_dma_0_mm_read_burstcount                       => read_dma_0_mm_read_burstcount,                     --                                              .burstcount
			read_dma_0_mm_read_byteenable                       => read_dma_0_mm_read_byteenable,                     --                                              .byteenable
			read_dma_0_mm_read_read                             => read_dma_0_mm_read_read,                           --                                              .read
			read_dma_0_mm_read_readdata                         => read_dma_0_mm_read_readdata,                       --                                              .readdata
			read_dma_0_mm_read_readdatavalid                    => read_dma_0_mm_read_readdatavalid,                  --                                              .readdatavalid
			video_dma_mm_read_address                           => video_dma_mm_read_address,                         --                             video_dma_mm_read.address
			video_dma_mm_read_waitrequest                       => video_dma_mm_read_waitrequest,                     --                                              .waitrequest
			video_dma_mm_read_burstcount                        => video_dma_mm_read_burstcount,                      --                                              .burstcount
			video_dma_mm_read_byteenable                        => video_dma_mm_read_byteenable,                      --                                              .byteenable
			video_dma_mm_read_read                              => video_dma_mm_read_read,                            --                                              .read
			video_dma_mm_read_readdata                          => video_dma_mm_read_readdata,                        --                                              .readdata
			video_dma_mm_read_readdatavalid                     => video_dma_mm_read_readdatavalid,                   --                                              .readdatavalid
			lpddr2_avl_1_address                                => mm_interconnect_1_lpddr2_avl_1_address,            --                                  lpddr2_avl_1.address
			lpddr2_avl_1_write                                  => mm_interconnect_1_lpddr2_avl_1_write,              --                                              .write
			lpddr2_avl_1_read                                   => mm_interconnect_1_lpddr2_avl_1_read,               --                                              .read
			lpddr2_avl_1_readdata                               => mm_interconnect_1_lpddr2_avl_1_readdata,           --                                              .readdata
			lpddr2_avl_1_writedata                              => mm_interconnect_1_lpddr2_avl_1_writedata,          --                                              .writedata
			lpddr2_avl_1_beginbursttransfer                     => mm_interconnect_1_lpddr2_avl_1_beginbursttransfer, --                                              .beginbursttransfer
			lpddr2_avl_1_burstcount                             => mm_interconnect_1_lpddr2_avl_1_burstcount,         --                                              .burstcount
			lpddr2_avl_1_byteenable                             => mm_interconnect_1_lpddr2_avl_1_byteenable,         --                                              .byteenable
			lpddr2_avl_1_readdatavalid                          => mm_interconnect_1_lpddr2_avl_1_readdatavalid,      --                                              .readdatavalid
			lpddr2_avl_1_waitrequest                            => mm_interconnect_1_lpddr2_avl_1_inv                 --                                              .waitrequest
		);

	mm_interconnect_2 : component HW_QSYS_mm_interconnect_2
		port map (
			clk_125_clk_clk                                     => clk_125_clk,                                       --                                   clk_125_clk.clk
			lpddr2_mp_cmd_reset_n_2_reset_bridge_in_reset_reset => rst_controller_004_reset_out_reset,                -- lpddr2_mp_cmd_reset_n_2_reset_bridge_in_reset.reset
			write_dma_0_reset_n_reset_bridge_in_reset_reset     => rst_controller_004_reset_out_reset,                --     write_dma_0_reset_n_reset_bridge_in_reset.reset
			write_dma_0_mm_write_address                        => write_dma_0_mm_write_address,                      --                          write_dma_0_mm_write.address
			write_dma_0_mm_write_waitrequest                    => write_dma_0_mm_write_waitrequest,                  --                                              .waitrequest
			write_dma_0_mm_write_burstcount                     => write_dma_0_mm_write_burstcount,                   --                                              .burstcount
			write_dma_0_mm_write_byteenable                     => write_dma_0_mm_write_byteenable,                   --                                              .byteenable
			write_dma_0_mm_write_write                          => write_dma_0_mm_write_write,                        --                                              .write
			write_dma_0_mm_write_writedata                      => write_dma_0_mm_write_writedata,                    --                                              .writedata
			lpddr2_avl_2_address                                => mm_interconnect_2_lpddr2_avl_2_address,            --                                  lpddr2_avl_2.address
			lpddr2_avl_2_write                                  => mm_interconnect_2_lpddr2_avl_2_write,              --                                              .write
			lpddr2_avl_2_read                                   => mm_interconnect_2_lpddr2_avl_2_read,               --                                              .read
			lpddr2_avl_2_readdata                               => mm_interconnect_2_lpddr2_avl_2_readdata,           --                                              .readdata
			lpddr2_avl_2_writedata                              => mm_interconnect_2_lpddr2_avl_2_writedata,          --                                              .writedata
			lpddr2_avl_2_beginbursttransfer                     => mm_interconnect_2_lpddr2_avl_2_beginbursttransfer, --                                              .beginbursttransfer
			lpddr2_avl_2_burstcount                             => mm_interconnect_2_lpddr2_avl_2_burstcount,         --                                              .burstcount
			lpddr2_avl_2_byteenable                             => mm_interconnect_2_lpddr2_avl_2_byteenable,         --                                              .byteenable
			lpddr2_avl_2_readdatavalid                          => mm_interconnect_2_lpddr2_avl_2_readdatavalid,      --                                              .readdatavalid
			lpddr2_avl_2_waitrequest                            => mm_interconnect_2_lpddr2_avl_2_inv                 --                                              .waitrequest
		);

	irq_mapper : component HW_QSYS_irq_mapper
		port map (
			clk           => clk_125_clk,                        --       clk.clk
			reset         => rst_controller_001_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,           -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,           -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,           -- receiver4.irq
			receiver5_irq => irq_mapper_receiver5_irq,           -- receiver5.irq
			receiver6_irq => irq_mapper_receiver6_irq,           -- receiver6.irq
			receiver7_irq => irq_mapper_receiver7_irq,           -- receiver7.irq
			receiver8_irq => irq_mapper_receiver8_irq,           -- receiver8.irq
			sender_irq    => cpu_0_irq_irq                       --    sender.irq
		);

	irq_mapper_001 : component HW_QSYS_irq_mapper_001
		port map (
			clk           => clk_125_clk,                        --       clk.clk
			reset         => rst_controller_002_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_001_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_001_receiver1_irq,       -- receiver1.irq
			sender_irq    => cpu_1_irq_irq                       --    sender.irq
		);

	irq_mapper_002 : component HW_QSYS_irq_mapper_001
		port map (
			clk           => clk_125_clk,                        --       clk.clk
			reset         => rst_controller_003_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_002_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_002_receiver1_irq,       -- receiver1.irq
			sender_irq    => cpu_2_irq_irq                       --    sender.irq
		);

	avalon_st_adapter : component HW_QSYS_avalon_st_adapter
		generic map (
			inBitsPerSymbol => 8,
			inUsePackets    => 1,
			inDataWidth     => 32,
			inChannelWidth  => 0,
			inErrorWidth    => 0,
			inUseEmptyPort  => 1,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 1,
			outDataWidth    => 32,
			outChannelWidth => 0,
			outErrorWidth   => 0,
			outUseEmptyPort => 1,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk        => video_pll_outclk0_clk,                 -- in_clk_0.clk
			in_rst_0_reset      => rst_controller_reset_out_reset,        -- in_rst_0.reset
			in_0_data           => video_fifo_out_data,                   --     in_0.data
			in_0_valid          => video_fifo_out_valid,                  --         .valid
			in_0_ready          => video_fifo_out_ready,                  --         .ready
			in_0_startofpacket  => video_fifo_out_startofpacket,          --         .startofpacket
			in_0_endofpacket    => video_fifo_out_endofpacket,            --         .endofpacket
			in_0_empty          => video_fifo_out_empty,                  --         .empty
			out_0_data          => avalon_st_adapter_out_0_data,          --    out_0.data
			out_0_valid         => avalon_st_adapter_out_0_valid,         --         .valid
			out_0_ready         => avalon_st_adapter_out_0_ready,         --         .ready
			out_0_startofpacket => avalon_st_adapter_out_0_startofpacket, --         .startofpacket
			out_0_endofpacket   => avalon_st_adapter_out_0_endofpacket,   --         .endofpacket
			out_0_empty         => avalon_st_adapter_out_0_empty          --         .empty
		);

	avalon_st_adapter_001 : component HW_QSYS_avalon_st_adapter_001
		generic map (
			inBitsPerSymbol => 8,
			inUsePackets    => 1,
			inDataWidth     => 32,
			inChannelWidth  => 0,
			inErrorWidth    => 0,
			inUseEmptyPort  => 1,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 0,
			outDataWidth    => 32,
			outChannelWidth => 0,
			outErrorWidth   => 0,
			outUseEmptyPort => 1,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 1
		)
		port map (
			in_clk_0_clk        => clk_125_clk,                               -- in_clk_0.clk
			in_rst_0_reset      => rst_controller_004_reset_out_reset,        -- in_rst_0.reset
			in_0_data           => video_dma_st_source_data,                  --     in_0.data
			in_0_valid          => video_dma_st_source_valid,                 --         .valid
			in_0_ready          => video_dma_st_source_ready,                 --         .ready
			in_0_startofpacket  => video_dma_st_source_startofpacket,         --         .startofpacket
			in_0_endofpacket    => video_dma_st_source_endofpacket,           --         .endofpacket
			in_0_empty          => video_dma_st_source_empty,                 --         .empty
			out_0_data          => avalon_st_adapter_001_out_0_data,          --    out_0.data
			out_0_valid         => avalon_st_adapter_001_out_0_valid,         --         .valid
			out_0_ready         => avalon_st_adapter_001_out_0_ready,         --         .ready
			out_0_startofpacket => avalon_st_adapter_001_out_0_startofpacket, --         .startofpacket
			out_0_endofpacket   => avalon_st_adapter_001_out_0_endofpacket,   --         .endofpacket
			out_0_empty         => avalon_st_adapter_001_out_0_empty          --         .empty
		);

	rst_controller : component HW_qsys_reset_controller_0
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_controller_0_reset_out_reset, -- reset_in0.reset
			clk            => video_pll_outclk0_clk,              --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component HW_qsys_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => cpu_0_debug_reset_request_reset,        -- reset_in0.reset
			reset_in1      => reset_controller_0_reset_out_reset,     -- reset_in1.reset
			clk            => clk_125_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_002 : component HW_qsys_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => cpu_1_debug_reset_request_reset,        -- reset_in0.reset
			reset_in1      => reset_controller_0_reset_out_reset,     -- reset_in1.reset
			clk            => clk_125_clk,                            --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_002_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_003 : component HW_qsys_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => cpu_2_debug_reset_request_reset,        -- reset_in0.reset
			reset_in1      => reset_controller_0_reset_out_reset,     -- reset_in1.reset
			clk            => clk_125_clk,                            --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_003_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_004 : component HW_qsys_reset_controller_0
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_controller_0_reset_out_reset, -- reset_in0.reset
			clk            => clk_125_clk,                        --       clk.clk
			reset_out      => rst_controller_004_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_005 : component HW_qsys_reset_controller_0
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_controller_0_reset_out_reset, -- reset_in0.reset
			clk            => clk_50_clk,                         --       clk.clk
			reset_out      => rst_controller_005_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	reset_controller_0_reset_out_reset_ports_inv <= not reset_controller_0_reset_out_reset;

	sd_cont_0_master_inv <= not mm_interconnect_0_sd_cont_0_master_waitrequest;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_lpddr2_avl_0_inv <= not lpddr2_avl_0_waitrequest;

	mm_interconnect_0_timer_0_s1_write_ports_inv <= not mm_interconnect_0_timer_0_s1_write;

	mm_interconnect_0_key_s1_write_ports_inv <= not mm_interconnect_0_key_s1_write;

	mm_interconnect_0_timer_1_s1_write_ports_inv <= not mm_interconnect_0_timer_1_s1_write;

	mm_interconnect_0_ledg_s1_write_ports_inv <= not mm_interconnect_0_ledg_s1_write;

	mm_interconnect_0_ledr_s1_write_ports_inv <= not mm_interconnect_0_ledr_s1_write;

	mm_interconnect_0_i2c_scl_s1_write_ports_inv <= not mm_interconnect_0_i2c_scl_s1_write;

	mm_interconnect_0_i2c_sda_s1_write_ports_inv <= not mm_interconnect_0_i2c_sda_s1_write;

	mm_interconnect_0_sd_cont_0_slave_inv <= not sd_cont_0_slave_waitrequest;

	mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_2_avalon_jtag_slave_write;

	mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write;

	mm_interconnect_1_lpddr2_avl_1_inv <= not lpddr2_avl_1_waitrequest;

	mm_interconnect_2_lpddr2_avl_2_inv <= not lpddr2_avl_2_waitrequest;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

	rst_controller_003_reset_out_reset_ports_inv <= not rst_controller_003_reset_out_reset;

	rst_controller_004_reset_out_reset_ports_inv <= not rst_controller_004_reset_out_reset;

	video_clk_clk <= video_pll_outclk0_clk;

end architecture rtl; -- of HW_QSYS
