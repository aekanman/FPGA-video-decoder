// HW_QSYS.v

// Generated using ACDS version 15.1 193

`timescale 1 ps / 1 ps
module HW_QSYS (
	);

	HW_QSYS_QSYS_0 qsys_0 (
	);

endmodule
